module Conwaylife(
  input          clock,
  input          reset,
  input          io_load,
  input  [255:0] io_data,
  output [255:0] io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg  regs_0_0; // @[Conwaylife.scala 10:17]
  reg  regs_0_1; // @[Conwaylife.scala 10:17]
  reg  regs_0_2; // @[Conwaylife.scala 10:17]
  reg  regs_0_3; // @[Conwaylife.scala 10:17]
  reg  regs_0_4; // @[Conwaylife.scala 10:17]
  reg  regs_0_5; // @[Conwaylife.scala 10:17]
  reg  regs_0_6; // @[Conwaylife.scala 10:17]
  reg  regs_0_7; // @[Conwaylife.scala 10:17]
  reg  regs_0_8; // @[Conwaylife.scala 10:17]
  reg  regs_0_9; // @[Conwaylife.scala 10:17]
  reg  regs_0_10; // @[Conwaylife.scala 10:17]
  reg  regs_0_11; // @[Conwaylife.scala 10:17]
  reg  regs_0_12; // @[Conwaylife.scala 10:17]
  reg  regs_0_13; // @[Conwaylife.scala 10:17]
  reg  regs_0_14; // @[Conwaylife.scala 10:17]
  reg  regs_0_15; // @[Conwaylife.scala 10:17]
  reg  regs_1_0; // @[Conwaylife.scala 10:17]
  reg  regs_1_1; // @[Conwaylife.scala 10:17]
  reg  regs_1_2; // @[Conwaylife.scala 10:17]
  reg  regs_1_3; // @[Conwaylife.scala 10:17]
  reg  regs_1_4; // @[Conwaylife.scala 10:17]
  reg  regs_1_5; // @[Conwaylife.scala 10:17]
  reg  regs_1_6; // @[Conwaylife.scala 10:17]
  reg  regs_1_7; // @[Conwaylife.scala 10:17]
  reg  regs_1_8; // @[Conwaylife.scala 10:17]
  reg  regs_1_9; // @[Conwaylife.scala 10:17]
  reg  regs_1_10; // @[Conwaylife.scala 10:17]
  reg  regs_1_11; // @[Conwaylife.scala 10:17]
  reg  regs_1_12; // @[Conwaylife.scala 10:17]
  reg  regs_1_13; // @[Conwaylife.scala 10:17]
  reg  regs_1_14; // @[Conwaylife.scala 10:17]
  reg  regs_1_15; // @[Conwaylife.scala 10:17]
  reg  regs_2_0; // @[Conwaylife.scala 10:17]
  reg  regs_2_1; // @[Conwaylife.scala 10:17]
  reg  regs_2_2; // @[Conwaylife.scala 10:17]
  reg  regs_2_3; // @[Conwaylife.scala 10:17]
  reg  regs_2_4; // @[Conwaylife.scala 10:17]
  reg  regs_2_5; // @[Conwaylife.scala 10:17]
  reg  regs_2_6; // @[Conwaylife.scala 10:17]
  reg  regs_2_7; // @[Conwaylife.scala 10:17]
  reg  regs_2_8; // @[Conwaylife.scala 10:17]
  reg  regs_2_9; // @[Conwaylife.scala 10:17]
  reg  regs_2_10; // @[Conwaylife.scala 10:17]
  reg  regs_2_11; // @[Conwaylife.scala 10:17]
  reg  regs_2_12; // @[Conwaylife.scala 10:17]
  reg  regs_2_13; // @[Conwaylife.scala 10:17]
  reg  regs_2_14; // @[Conwaylife.scala 10:17]
  reg  regs_2_15; // @[Conwaylife.scala 10:17]
  reg  regs_3_0; // @[Conwaylife.scala 10:17]
  reg  regs_3_1; // @[Conwaylife.scala 10:17]
  reg  regs_3_2; // @[Conwaylife.scala 10:17]
  reg  regs_3_3; // @[Conwaylife.scala 10:17]
  reg  regs_3_4; // @[Conwaylife.scala 10:17]
  reg  regs_3_5; // @[Conwaylife.scala 10:17]
  reg  regs_3_6; // @[Conwaylife.scala 10:17]
  reg  regs_3_7; // @[Conwaylife.scala 10:17]
  reg  regs_3_8; // @[Conwaylife.scala 10:17]
  reg  regs_3_9; // @[Conwaylife.scala 10:17]
  reg  regs_3_10; // @[Conwaylife.scala 10:17]
  reg  regs_3_11; // @[Conwaylife.scala 10:17]
  reg  regs_3_12; // @[Conwaylife.scala 10:17]
  reg  regs_3_13; // @[Conwaylife.scala 10:17]
  reg  regs_3_14; // @[Conwaylife.scala 10:17]
  reg  regs_3_15; // @[Conwaylife.scala 10:17]
  reg  regs_4_0; // @[Conwaylife.scala 10:17]
  reg  regs_4_1; // @[Conwaylife.scala 10:17]
  reg  regs_4_2; // @[Conwaylife.scala 10:17]
  reg  regs_4_3; // @[Conwaylife.scala 10:17]
  reg  regs_4_4; // @[Conwaylife.scala 10:17]
  reg  regs_4_5; // @[Conwaylife.scala 10:17]
  reg  regs_4_6; // @[Conwaylife.scala 10:17]
  reg  regs_4_7; // @[Conwaylife.scala 10:17]
  reg  regs_4_8; // @[Conwaylife.scala 10:17]
  reg  regs_4_9; // @[Conwaylife.scala 10:17]
  reg  regs_4_10; // @[Conwaylife.scala 10:17]
  reg  regs_4_11; // @[Conwaylife.scala 10:17]
  reg  regs_4_12; // @[Conwaylife.scala 10:17]
  reg  regs_4_13; // @[Conwaylife.scala 10:17]
  reg  regs_4_14; // @[Conwaylife.scala 10:17]
  reg  regs_4_15; // @[Conwaylife.scala 10:17]
  reg  regs_5_0; // @[Conwaylife.scala 10:17]
  reg  regs_5_1; // @[Conwaylife.scala 10:17]
  reg  regs_5_2; // @[Conwaylife.scala 10:17]
  reg  regs_5_3; // @[Conwaylife.scala 10:17]
  reg  regs_5_4; // @[Conwaylife.scala 10:17]
  reg  regs_5_5; // @[Conwaylife.scala 10:17]
  reg  regs_5_6; // @[Conwaylife.scala 10:17]
  reg  regs_5_7; // @[Conwaylife.scala 10:17]
  reg  regs_5_8; // @[Conwaylife.scala 10:17]
  reg  regs_5_9; // @[Conwaylife.scala 10:17]
  reg  regs_5_10; // @[Conwaylife.scala 10:17]
  reg  regs_5_11; // @[Conwaylife.scala 10:17]
  reg  regs_5_12; // @[Conwaylife.scala 10:17]
  reg  regs_5_13; // @[Conwaylife.scala 10:17]
  reg  regs_5_14; // @[Conwaylife.scala 10:17]
  reg  regs_5_15; // @[Conwaylife.scala 10:17]
  reg  regs_6_0; // @[Conwaylife.scala 10:17]
  reg  regs_6_1; // @[Conwaylife.scala 10:17]
  reg  regs_6_2; // @[Conwaylife.scala 10:17]
  reg  regs_6_3; // @[Conwaylife.scala 10:17]
  reg  regs_6_4; // @[Conwaylife.scala 10:17]
  reg  regs_6_5; // @[Conwaylife.scala 10:17]
  reg  regs_6_6; // @[Conwaylife.scala 10:17]
  reg  regs_6_7; // @[Conwaylife.scala 10:17]
  reg  regs_6_8; // @[Conwaylife.scala 10:17]
  reg  regs_6_9; // @[Conwaylife.scala 10:17]
  reg  regs_6_10; // @[Conwaylife.scala 10:17]
  reg  regs_6_11; // @[Conwaylife.scala 10:17]
  reg  regs_6_12; // @[Conwaylife.scala 10:17]
  reg  regs_6_13; // @[Conwaylife.scala 10:17]
  reg  regs_6_14; // @[Conwaylife.scala 10:17]
  reg  regs_6_15; // @[Conwaylife.scala 10:17]
  reg  regs_7_0; // @[Conwaylife.scala 10:17]
  reg  regs_7_1; // @[Conwaylife.scala 10:17]
  reg  regs_7_2; // @[Conwaylife.scala 10:17]
  reg  regs_7_3; // @[Conwaylife.scala 10:17]
  reg  regs_7_4; // @[Conwaylife.scala 10:17]
  reg  regs_7_5; // @[Conwaylife.scala 10:17]
  reg  regs_7_6; // @[Conwaylife.scala 10:17]
  reg  regs_7_7; // @[Conwaylife.scala 10:17]
  reg  regs_7_8; // @[Conwaylife.scala 10:17]
  reg  regs_7_9; // @[Conwaylife.scala 10:17]
  reg  regs_7_10; // @[Conwaylife.scala 10:17]
  reg  regs_7_11; // @[Conwaylife.scala 10:17]
  reg  regs_7_12; // @[Conwaylife.scala 10:17]
  reg  regs_7_13; // @[Conwaylife.scala 10:17]
  reg  regs_7_14; // @[Conwaylife.scala 10:17]
  reg  regs_7_15; // @[Conwaylife.scala 10:17]
  reg  regs_8_0; // @[Conwaylife.scala 10:17]
  reg  regs_8_1; // @[Conwaylife.scala 10:17]
  reg  regs_8_2; // @[Conwaylife.scala 10:17]
  reg  regs_8_3; // @[Conwaylife.scala 10:17]
  reg  regs_8_4; // @[Conwaylife.scala 10:17]
  reg  regs_8_5; // @[Conwaylife.scala 10:17]
  reg  regs_8_6; // @[Conwaylife.scala 10:17]
  reg  regs_8_7; // @[Conwaylife.scala 10:17]
  reg  regs_8_8; // @[Conwaylife.scala 10:17]
  reg  regs_8_9; // @[Conwaylife.scala 10:17]
  reg  regs_8_10; // @[Conwaylife.scala 10:17]
  reg  regs_8_11; // @[Conwaylife.scala 10:17]
  reg  regs_8_12; // @[Conwaylife.scala 10:17]
  reg  regs_8_13; // @[Conwaylife.scala 10:17]
  reg  regs_8_14; // @[Conwaylife.scala 10:17]
  reg  regs_8_15; // @[Conwaylife.scala 10:17]
  reg  regs_9_0; // @[Conwaylife.scala 10:17]
  reg  regs_9_1; // @[Conwaylife.scala 10:17]
  reg  regs_9_2; // @[Conwaylife.scala 10:17]
  reg  regs_9_3; // @[Conwaylife.scala 10:17]
  reg  regs_9_4; // @[Conwaylife.scala 10:17]
  reg  regs_9_5; // @[Conwaylife.scala 10:17]
  reg  regs_9_6; // @[Conwaylife.scala 10:17]
  reg  regs_9_7; // @[Conwaylife.scala 10:17]
  reg  regs_9_8; // @[Conwaylife.scala 10:17]
  reg  regs_9_9; // @[Conwaylife.scala 10:17]
  reg  regs_9_10; // @[Conwaylife.scala 10:17]
  reg  regs_9_11; // @[Conwaylife.scala 10:17]
  reg  regs_9_12; // @[Conwaylife.scala 10:17]
  reg  regs_9_13; // @[Conwaylife.scala 10:17]
  reg  regs_9_14; // @[Conwaylife.scala 10:17]
  reg  regs_9_15; // @[Conwaylife.scala 10:17]
  reg  regs_10_0; // @[Conwaylife.scala 10:17]
  reg  regs_10_1; // @[Conwaylife.scala 10:17]
  reg  regs_10_2; // @[Conwaylife.scala 10:17]
  reg  regs_10_3; // @[Conwaylife.scala 10:17]
  reg  regs_10_4; // @[Conwaylife.scala 10:17]
  reg  regs_10_5; // @[Conwaylife.scala 10:17]
  reg  regs_10_6; // @[Conwaylife.scala 10:17]
  reg  regs_10_7; // @[Conwaylife.scala 10:17]
  reg  regs_10_8; // @[Conwaylife.scala 10:17]
  reg  regs_10_9; // @[Conwaylife.scala 10:17]
  reg  regs_10_10; // @[Conwaylife.scala 10:17]
  reg  regs_10_11; // @[Conwaylife.scala 10:17]
  reg  regs_10_12; // @[Conwaylife.scala 10:17]
  reg  regs_10_13; // @[Conwaylife.scala 10:17]
  reg  regs_10_14; // @[Conwaylife.scala 10:17]
  reg  regs_10_15; // @[Conwaylife.scala 10:17]
  reg  regs_11_0; // @[Conwaylife.scala 10:17]
  reg  regs_11_1; // @[Conwaylife.scala 10:17]
  reg  regs_11_2; // @[Conwaylife.scala 10:17]
  reg  regs_11_3; // @[Conwaylife.scala 10:17]
  reg  regs_11_4; // @[Conwaylife.scala 10:17]
  reg  regs_11_5; // @[Conwaylife.scala 10:17]
  reg  regs_11_6; // @[Conwaylife.scala 10:17]
  reg  regs_11_7; // @[Conwaylife.scala 10:17]
  reg  regs_11_8; // @[Conwaylife.scala 10:17]
  reg  regs_11_9; // @[Conwaylife.scala 10:17]
  reg  regs_11_10; // @[Conwaylife.scala 10:17]
  reg  regs_11_11; // @[Conwaylife.scala 10:17]
  reg  regs_11_12; // @[Conwaylife.scala 10:17]
  reg  regs_11_13; // @[Conwaylife.scala 10:17]
  reg  regs_11_14; // @[Conwaylife.scala 10:17]
  reg  regs_11_15; // @[Conwaylife.scala 10:17]
  reg  regs_12_0; // @[Conwaylife.scala 10:17]
  reg  regs_12_1; // @[Conwaylife.scala 10:17]
  reg  regs_12_2; // @[Conwaylife.scala 10:17]
  reg  regs_12_3; // @[Conwaylife.scala 10:17]
  reg  regs_12_4; // @[Conwaylife.scala 10:17]
  reg  regs_12_5; // @[Conwaylife.scala 10:17]
  reg  regs_12_6; // @[Conwaylife.scala 10:17]
  reg  regs_12_7; // @[Conwaylife.scala 10:17]
  reg  regs_12_8; // @[Conwaylife.scala 10:17]
  reg  regs_12_9; // @[Conwaylife.scala 10:17]
  reg  regs_12_10; // @[Conwaylife.scala 10:17]
  reg  regs_12_11; // @[Conwaylife.scala 10:17]
  reg  regs_12_12; // @[Conwaylife.scala 10:17]
  reg  regs_12_13; // @[Conwaylife.scala 10:17]
  reg  regs_12_14; // @[Conwaylife.scala 10:17]
  reg  regs_12_15; // @[Conwaylife.scala 10:17]
  reg  regs_13_0; // @[Conwaylife.scala 10:17]
  reg  regs_13_1; // @[Conwaylife.scala 10:17]
  reg  regs_13_2; // @[Conwaylife.scala 10:17]
  reg  regs_13_3; // @[Conwaylife.scala 10:17]
  reg  regs_13_4; // @[Conwaylife.scala 10:17]
  reg  regs_13_5; // @[Conwaylife.scala 10:17]
  reg  regs_13_6; // @[Conwaylife.scala 10:17]
  reg  regs_13_7; // @[Conwaylife.scala 10:17]
  reg  regs_13_8; // @[Conwaylife.scala 10:17]
  reg  regs_13_9; // @[Conwaylife.scala 10:17]
  reg  regs_13_10; // @[Conwaylife.scala 10:17]
  reg  regs_13_11; // @[Conwaylife.scala 10:17]
  reg  regs_13_12; // @[Conwaylife.scala 10:17]
  reg  regs_13_13; // @[Conwaylife.scala 10:17]
  reg  regs_13_14; // @[Conwaylife.scala 10:17]
  reg  regs_13_15; // @[Conwaylife.scala 10:17]
  reg  regs_14_0; // @[Conwaylife.scala 10:17]
  reg  regs_14_1; // @[Conwaylife.scala 10:17]
  reg  regs_14_2; // @[Conwaylife.scala 10:17]
  reg  regs_14_3; // @[Conwaylife.scala 10:17]
  reg  regs_14_4; // @[Conwaylife.scala 10:17]
  reg  regs_14_5; // @[Conwaylife.scala 10:17]
  reg  regs_14_6; // @[Conwaylife.scala 10:17]
  reg  regs_14_7; // @[Conwaylife.scala 10:17]
  reg  regs_14_8; // @[Conwaylife.scala 10:17]
  reg  regs_14_9; // @[Conwaylife.scala 10:17]
  reg  regs_14_10; // @[Conwaylife.scala 10:17]
  reg  regs_14_11; // @[Conwaylife.scala 10:17]
  reg  regs_14_12; // @[Conwaylife.scala 10:17]
  reg  regs_14_13; // @[Conwaylife.scala 10:17]
  reg  regs_14_14; // @[Conwaylife.scala 10:17]
  reg  regs_14_15; // @[Conwaylife.scala 10:17]
  reg  regs_15_0; // @[Conwaylife.scala 10:17]
  reg  regs_15_1; // @[Conwaylife.scala 10:17]
  reg  regs_15_2; // @[Conwaylife.scala 10:17]
  reg  regs_15_3; // @[Conwaylife.scala 10:17]
  reg  regs_15_4; // @[Conwaylife.scala 10:17]
  reg  regs_15_5; // @[Conwaylife.scala 10:17]
  reg  regs_15_6; // @[Conwaylife.scala 10:17]
  reg  regs_15_7; // @[Conwaylife.scala 10:17]
  reg  regs_15_8; // @[Conwaylife.scala 10:17]
  reg  regs_15_9; // @[Conwaylife.scala 10:17]
  reg  regs_15_10; // @[Conwaylife.scala 10:17]
  reg  regs_15_11; // @[Conwaylife.scala 10:17]
  reg  regs_15_12; // @[Conwaylife.scala 10:17]
  reg  regs_15_13; // @[Conwaylife.scala 10:17]
  reg  regs_15_14; // @[Conwaylife.scala 10:17]
  reg  regs_15_15; // @[Conwaylife.scala 10:17]
  wire [1:0] _T_256 = regs_15_15 + regs_15_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1024 = {{1'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_257 = _T_256 + _GEN_1024; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1025 = {{2'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_258 = _T_257 + _GEN_1025; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1026 = {{3'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_259 = _T_258 + _GEN_1026; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1027 = {{4'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_260 = _T_259 + _GEN_1027; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1028 = {{5'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_261 = _T_260 + _GEN_1028; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1029 = {{6'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_262 = _T_261 + _GEN_1029; // @[Conwaylife.scala 31:34]
  wire  _T_263 = _T_262 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_264 = _T_262 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_265 = _T_262 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_266 = regs_15_0 + regs_15_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1030 = {{1'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_267 = _T_266 + _GEN_1030; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1031 = {{2'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_268 = _T_267 + _GEN_1031; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1032 = {{3'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_269 = _T_268 + _GEN_1032; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1033 = {{4'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_270 = _T_269 + _GEN_1033; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1034 = {{5'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_271 = _T_270 + _GEN_1034; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1035 = {{6'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_272 = _T_271 + _GEN_1035; // @[Conwaylife.scala 31:34]
  wire  _T_273 = _T_272 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_274 = _T_272 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_275 = _T_272 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_276 = regs_15_1 + regs_15_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1036 = {{1'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_277 = _T_276 + _GEN_1036; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1037 = {{2'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_278 = _T_277 + _GEN_1037; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1038 = {{3'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_279 = _T_278 + _GEN_1038; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1039 = {{4'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_280 = _T_279 + _GEN_1039; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1040 = {{5'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_281 = _T_280 + _GEN_1040; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1041 = {{6'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_282 = _T_281 + _GEN_1041; // @[Conwaylife.scala 31:34]
  wire  _T_283 = _T_282 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_284 = _T_282 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_285 = _T_282 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_286 = regs_15_2 + regs_15_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1042 = {{1'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_287 = _T_286 + _GEN_1042; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1043 = {{2'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_288 = _T_287 + _GEN_1043; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1044 = {{3'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_289 = _T_288 + _GEN_1044; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1045 = {{4'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_290 = _T_289 + _GEN_1045; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1046 = {{5'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_291 = _T_290 + _GEN_1046; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1047 = {{6'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_292 = _T_291 + _GEN_1047; // @[Conwaylife.scala 31:34]
  wire  _T_293 = _T_292 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_294 = _T_292 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_295 = _T_292 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_296 = regs_15_3 + regs_15_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1048 = {{1'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_297 = _T_296 + _GEN_1048; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1049 = {{2'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_298 = _T_297 + _GEN_1049; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1050 = {{3'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_299 = _T_298 + _GEN_1050; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1051 = {{4'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_300 = _T_299 + _GEN_1051; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1052 = {{5'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_301 = _T_300 + _GEN_1052; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1053 = {{6'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_302 = _T_301 + _GEN_1053; // @[Conwaylife.scala 31:34]
  wire  _T_303 = _T_302 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_304 = _T_302 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_305 = _T_302 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_306 = regs_15_4 + regs_15_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1054 = {{1'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_307 = _T_306 + _GEN_1054; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1055 = {{2'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_308 = _T_307 + _GEN_1055; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1056 = {{3'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_309 = _T_308 + _GEN_1056; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1057 = {{4'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_310 = _T_309 + _GEN_1057; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1058 = {{5'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_311 = _T_310 + _GEN_1058; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1059 = {{6'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_312 = _T_311 + _GEN_1059; // @[Conwaylife.scala 31:34]
  wire  _T_313 = _T_312 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_314 = _T_312 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_315 = _T_312 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_316 = regs_15_5 + regs_15_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1060 = {{1'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_317 = _T_316 + _GEN_1060; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1061 = {{2'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_318 = _T_317 + _GEN_1061; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1062 = {{3'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_319 = _T_318 + _GEN_1062; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1063 = {{4'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_320 = _T_319 + _GEN_1063; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1064 = {{5'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_321 = _T_320 + _GEN_1064; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1065 = {{6'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_322 = _T_321 + _GEN_1065; // @[Conwaylife.scala 31:34]
  wire  _T_323 = _T_322 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_324 = _T_322 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_325 = _T_322 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_326 = regs_15_6 + regs_15_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1066 = {{1'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_327 = _T_326 + _GEN_1066; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1067 = {{2'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_328 = _T_327 + _GEN_1067; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1068 = {{3'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_329 = _T_328 + _GEN_1068; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1069 = {{4'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_330 = _T_329 + _GEN_1069; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1070 = {{5'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_331 = _T_330 + _GEN_1070; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1071 = {{6'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_332 = _T_331 + _GEN_1071; // @[Conwaylife.scala 31:34]
  wire  _T_333 = _T_332 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_334 = _T_332 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_335 = _T_332 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_336 = regs_15_7 + regs_15_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1072 = {{1'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_337 = _T_336 + _GEN_1072; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1073 = {{2'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_338 = _T_337 + _GEN_1073; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1074 = {{3'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_339 = _T_338 + _GEN_1074; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1075 = {{4'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_340 = _T_339 + _GEN_1075; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1076 = {{5'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_341 = _T_340 + _GEN_1076; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1077 = {{6'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_342 = _T_341 + _GEN_1077; // @[Conwaylife.scala 31:34]
  wire  _T_343 = _T_342 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_344 = _T_342 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_345 = _T_342 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_346 = regs_15_8 + regs_15_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1078 = {{1'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_347 = _T_346 + _GEN_1078; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1079 = {{2'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_348 = _T_347 + _GEN_1079; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1080 = {{3'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_349 = _T_348 + _GEN_1080; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1081 = {{4'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_350 = _T_349 + _GEN_1081; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1082 = {{5'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_351 = _T_350 + _GEN_1082; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1083 = {{6'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_352 = _T_351 + _GEN_1083; // @[Conwaylife.scala 31:34]
  wire  _T_353 = _T_352 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_354 = _T_352 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_355 = _T_352 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_356 = regs_15_9 + regs_15_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1084 = {{1'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_357 = _T_356 + _GEN_1084; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1085 = {{2'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_358 = _T_357 + _GEN_1085; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1086 = {{3'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_359 = _T_358 + _GEN_1086; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1087 = {{4'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_360 = _T_359 + _GEN_1087; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1088 = {{5'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_361 = _T_360 + _GEN_1088; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1089 = {{6'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_362 = _T_361 + _GEN_1089; // @[Conwaylife.scala 31:34]
  wire  _T_363 = _T_362 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_364 = _T_362 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_365 = _T_362 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_366 = regs_15_10 + regs_15_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1090 = {{1'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_367 = _T_366 + _GEN_1090; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1091 = {{2'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_368 = _T_367 + _GEN_1091; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1092 = {{3'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_369 = _T_368 + _GEN_1092; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1093 = {{4'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_370 = _T_369 + _GEN_1093; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1094 = {{5'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_371 = _T_370 + _GEN_1094; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1095 = {{6'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_372 = _T_371 + _GEN_1095; // @[Conwaylife.scala 31:34]
  wire  _T_373 = _T_372 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_374 = _T_372 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_375 = _T_372 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_376 = regs_15_11 + regs_15_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1096 = {{1'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_377 = _T_376 + _GEN_1096; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1097 = {{2'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_378 = _T_377 + _GEN_1097; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1098 = {{3'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_379 = _T_378 + _GEN_1098; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1099 = {{4'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_380 = _T_379 + _GEN_1099; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1100 = {{5'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_381 = _T_380 + _GEN_1100; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1101 = {{6'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_382 = _T_381 + _GEN_1101; // @[Conwaylife.scala 31:34]
  wire  _T_383 = _T_382 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_384 = _T_382 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_385 = _T_382 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_386 = regs_15_12 + regs_15_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1102 = {{1'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_387 = _T_386 + _GEN_1102; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1103 = {{2'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_388 = _T_387 + _GEN_1103; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1104 = {{3'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_389 = _T_388 + _GEN_1104; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1105 = {{4'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_390 = _T_389 + _GEN_1105; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1106 = {{5'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_391 = _T_390 + _GEN_1106; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1107 = {{6'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_392 = _T_391 + _GEN_1107; // @[Conwaylife.scala 31:34]
  wire  _T_393 = _T_392 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_394 = _T_392 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_395 = _T_392 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_396 = regs_15_13 + regs_15_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1108 = {{1'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_397 = _T_396 + _GEN_1108; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1109 = {{2'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_398 = _T_397 + _GEN_1109; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1110 = {{3'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_399 = _T_398 + _GEN_1110; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1111 = {{4'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_400 = _T_399 + _GEN_1111; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1112 = {{5'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_401 = _T_400 + _GEN_1112; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1113 = {{6'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_402 = _T_401 + _GEN_1113; // @[Conwaylife.scala 31:34]
  wire  _T_403 = _T_402 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_404 = _T_402 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_405 = _T_402 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_406 = regs_15_14 + regs_15_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1114 = {{1'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_407 = _T_406 + _GEN_1114; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1115 = {{2'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_408 = _T_407 + _GEN_1115; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1116 = {{3'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_409 = _T_408 + _GEN_1116; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1117 = {{4'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_410 = _T_409 + _GEN_1117; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1118 = {{5'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_411 = _T_410 + _GEN_1118; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1119 = {{6'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_412 = _T_411 + _GEN_1119; // @[Conwaylife.scala 31:34]
  wire  _T_413 = _T_412 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_414 = _T_412 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_415 = _T_412 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_416 = regs_0_15 + regs_0_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1120 = {{1'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_417 = _T_416 + _GEN_1120; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1121 = {{2'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_418 = _T_417 + _GEN_1121; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1122 = {{3'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_419 = _T_418 + _GEN_1122; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1123 = {{4'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_420 = _T_419 + _GEN_1123; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1124 = {{5'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_421 = _T_420 + _GEN_1124; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1125 = {{6'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_422 = _T_421 + _GEN_1125; // @[Conwaylife.scala 31:34]
  wire  _T_423 = _T_422 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_424 = _T_422 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_425 = _T_422 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_426 = regs_0_0 + regs_0_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1126 = {{1'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_427 = _T_426 + _GEN_1126; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1127 = {{2'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_428 = _T_427 + _GEN_1127; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1128 = {{3'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_429 = _T_428 + _GEN_1128; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1129 = {{4'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_430 = _T_429 + _GEN_1129; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1130 = {{5'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_431 = _T_430 + _GEN_1130; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1131 = {{6'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_432 = _T_431 + _GEN_1131; // @[Conwaylife.scala 31:34]
  wire  _T_433 = _T_432 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_434 = _T_432 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_435 = _T_432 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_436 = regs_0_1 + regs_0_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1132 = {{1'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_437 = _T_436 + _GEN_1132; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1133 = {{2'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_438 = _T_437 + _GEN_1133; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1134 = {{3'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_439 = _T_438 + _GEN_1134; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1135 = {{4'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_440 = _T_439 + _GEN_1135; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1136 = {{5'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_441 = _T_440 + _GEN_1136; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1137 = {{6'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_442 = _T_441 + _GEN_1137; // @[Conwaylife.scala 31:34]
  wire  _T_443 = _T_442 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_444 = _T_442 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_445 = _T_442 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_446 = regs_0_2 + regs_0_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1138 = {{1'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_447 = _T_446 + _GEN_1138; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1139 = {{2'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_448 = _T_447 + _GEN_1139; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1140 = {{3'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_449 = _T_448 + _GEN_1140; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1141 = {{4'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_450 = _T_449 + _GEN_1141; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1142 = {{5'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_451 = _T_450 + _GEN_1142; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1143 = {{6'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_452 = _T_451 + _GEN_1143; // @[Conwaylife.scala 31:34]
  wire  _T_453 = _T_452 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_454 = _T_452 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_455 = _T_452 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_456 = regs_0_3 + regs_0_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1144 = {{1'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_457 = _T_456 + _GEN_1144; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1145 = {{2'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_458 = _T_457 + _GEN_1145; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1146 = {{3'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_459 = _T_458 + _GEN_1146; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1147 = {{4'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_460 = _T_459 + _GEN_1147; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1148 = {{5'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_461 = _T_460 + _GEN_1148; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1149 = {{6'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_462 = _T_461 + _GEN_1149; // @[Conwaylife.scala 31:34]
  wire  _T_463 = _T_462 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_464 = _T_462 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_465 = _T_462 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_466 = regs_0_4 + regs_0_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1150 = {{1'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_467 = _T_466 + _GEN_1150; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1151 = {{2'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_468 = _T_467 + _GEN_1151; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1152 = {{3'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_469 = _T_468 + _GEN_1152; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1153 = {{4'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_470 = _T_469 + _GEN_1153; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1154 = {{5'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_471 = _T_470 + _GEN_1154; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1155 = {{6'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_472 = _T_471 + _GEN_1155; // @[Conwaylife.scala 31:34]
  wire  _T_473 = _T_472 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_474 = _T_472 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_475 = _T_472 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_476 = regs_0_5 + regs_0_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1156 = {{1'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_477 = _T_476 + _GEN_1156; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1157 = {{2'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_478 = _T_477 + _GEN_1157; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1158 = {{3'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_479 = _T_478 + _GEN_1158; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1159 = {{4'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_480 = _T_479 + _GEN_1159; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1160 = {{5'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_481 = _T_480 + _GEN_1160; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1161 = {{6'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_482 = _T_481 + _GEN_1161; // @[Conwaylife.scala 31:34]
  wire  _T_483 = _T_482 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_484 = _T_482 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_485 = _T_482 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_486 = regs_0_6 + regs_0_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1162 = {{1'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_487 = _T_486 + _GEN_1162; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1163 = {{2'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_488 = _T_487 + _GEN_1163; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1164 = {{3'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_489 = _T_488 + _GEN_1164; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1165 = {{4'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_490 = _T_489 + _GEN_1165; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1166 = {{5'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_491 = _T_490 + _GEN_1166; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1167 = {{6'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_492 = _T_491 + _GEN_1167; // @[Conwaylife.scala 31:34]
  wire  _T_493 = _T_492 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_494 = _T_492 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_495 = _T_492 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_496 = regs_0_7 + regs_0_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1168 = {{1'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_497 = _T_496 + _GEN_1168; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1169 = {{2'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_498 = _T_497 + _GEN_1169; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1170 = {{3'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_499 = _T_498 + _GEN_1170; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1171 = {{4'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_500 = _T_499 + _GEN_1171; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1172 = {{5'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_501 = _T_500 + _GEN_1172; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1173 = {{6'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_502 = _T_501 + _GEN_1173; // @[Conwaylife.scala 31:34]
  wire  _T_503 = _T_502 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_504 = _T_502 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_505 = _T_502 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_506 = regs_0_8 + regs_0_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1174 = {{1'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_507 = _T_506 + _GEN_1174; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1175 = {{2'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_508 = _T_507 + _GEN_1175; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1176 = {{3'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_509 = _T_508 + _GEN_1176; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1177 = {{4'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_510 = _T_509 + _GEN_1177; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1178 = {{5'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_511 = _T_510 + _GEN_1178; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1179 = {{6'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_512 = _T_511 + _GEN_1179; // @[Conwaylife.scala 31:34]
  wire  _T_513 = _T_512 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_514 = _T_512 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_515 = _T_512 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_516 = regs_0_9 + regs_0_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1180 = {{1'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_517 = _T_516 + _GEN_1180; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1181 = {{2'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_518 = _T_517 + _GEN_1181; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1182 = {{3'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_519 = _T_518 + _GEN_1182; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1183 = {{4'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_520 = _T_519 + _GEN_1183; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1184 = {{5'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_521 = _T_520 + _GEN_1184; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1185 = {{6'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_522 = _T_521 + _GEN_1185; // @[Conwaylife.scala 31:34]
  wire  _T_523 = _T_522 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_524 = _T_522 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_525 = _T_522 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_526 = regs_0_10 + regs_0_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1186 = {{1'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_527 = _T_526 + _GEN_1186; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1187 = {{2'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_528 = _T_527 + _GEN_1187; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1188 = {{3'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_529 = _T_528 + _GEN_1188; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1189 = {{4'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_530 = _T_529 + _GEN_1189; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1190 = {{5'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_531 = _T_530 + _GEN_1190; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1191 = {{6'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_532 = _T_531 + _GEN_1191; // @[Conwaylife.scala 31:34]
  wire  _T_533 = _T_532 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_534 = _T_532 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_535 = _T_532 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_536 = regs_0_11 + regs_0_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1192 = {{1'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_537 = _T_536 + _GEN_1192; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1193 = {{2'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_538 = _T_537 + _GEN_1193; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1194 = {{3'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_539 = _T_538 + _GEN_1194; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1195 = {{4'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_540 = _T_539 + _GEN_1195; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1196 = {{5'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_541 = _T_540 + _GEN_1196; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1197 = {{6'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_542 = _T_541 + _GEN_1197; // @[Conwaylife.scala 31:34]
  wire  _T_543 = _T_542 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_544 = _T_542 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_545 = _T_542 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_546 = regs_0_12 + regs_0_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1198 = {{1'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_547 = _T_546 + _GEN_1198; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1199 = {{2'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_548 = _T_547 + _GEN_1199; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1200 = {{3'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_549 = _T_548 + _GEN_1200; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1201 = {{4'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_550 = _T_549 + _GEN_1201; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1202 = {{5'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_551 = _T_550 + _GEN_1202; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1203 = {{6'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_552 = _T_551 + _GEN_1203; // @[Conwaylife.scala 31:34]
  wire  _T_553 = _T_552 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_554 = _T_552 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_555 = _T_552 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_556 = regs_0_13 + regs_0_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1204 = {{1'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_557 = _T_556 + _GEN_1204; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1205 = {{2'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_558 = _T_557 + _GEN_1205; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1206 = {{3'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_559 = _T_558 + _GEN_1206; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1207 = {{4'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_560 = _T_559 + _GEN_1207; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1208 = {{5'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_561 = _T_560 + _GEN_1208; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1209 = {{6'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_562 = _T_561 + _GEN_1209; // @[Conwaylife.scala 31:34]
  wire  _T_563 = _T_562 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_564 = _T_562 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_565 = _T_562 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_566 = regs_0_14 + regs_0_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1210 = {{1'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_567 = _T_566 + _GEN_1210; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1211 = {{2'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_568 = _T_567 + _GEN_1211; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1212 = {{3'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_569 = _T_568 + _GEN_1212; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1213 = {{4'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_570 = _T_569 + _GEN_1213; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1214 = {{5'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_571 = _T_570 + _GEN_1214; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1215 = {{6'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_572 = _T_571 + _GEN_1215; // @[Conwaylife.scala 31:34]
  wire  _T_573 = _T_572 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_574 = _T_572 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_575 = _T_572 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_576 = regs_1_15 + regs_1_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1216 = {{1'd0}, regs_1_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_577 = _T_576 + _GEN_1216; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1217 = {{2'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_578 = _T_577 + _GEN_1217; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1218 = {{3'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_579 = _T_578 + _GEN_1218; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1219 = {{4'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_580 = _T_579 + _GEN_1219; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1220 = {{5'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_581 = _T_580 + _GEN_1220; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1221 = {{6'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_582 = _T_581 + _GEN_1221; // @[Conwaylife.scala 31:34]
  wire  _T_583 = _T_582 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_584 = _T_582 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_585 = _T_582 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_586 = regs_1_0 + regs_1_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1222 = {{1'd0}, regs_1_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_587 = _T_586 + _GEN_1222; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1223 = {{2'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_588 = _T_587 + _GEN_1223; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1224 = {{3'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_589 = _T_588 + _GEN_1224; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1225 = {{4'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_590 = _T_589 + _GEN_1225; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1226 = {{5'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_591 = _T_590 + _GEN_1226; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1227 = {{6'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_592 = _T_591 + _GEN_1227; // @[Conwaylife.scala 31:34]
  wire  _T_593 = _T_592 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_594 = _T_592 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_595 = _T_592 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_596 = regs_1_1 + regs_1_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1228 = {{1'd0}, regs_1_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_597 = _T_596 + _GEN_1228; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1229 = {{2'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_598 = _T_597 + _GEN_1229; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1230 = {{3'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_599 = _T_598 + _GEN_1230; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1231 = {{4'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_600 = _T_599 + _GEN_1231; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1232 = {{5'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_601 = _T_600 + _GEN_1232; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1233 = {{6'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_602 = _T_601 + _GEN_1233; // @[Conwaylife.scala 31:34]
  wire  _T_603 = _T_602 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_604 = _T_602 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_605 = _T_602 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_606 = regs_1_2 + regs_1_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1234 = {{1'd0}, regs_1_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_607 = _T_606 + _GEN_1234; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1235 = {{2'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_608 = _T_607 + _GEN_1235; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1236 = {{3'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_609 = _T_608 + _GEN_1236; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1237 = {{4'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_610 = _T_609 + _GEN_1237; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1238 = {{5'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_611 = _T_610 + _GEN_1238; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1239 = {{6'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_612 = _T_611 + _GEN_1239; // @[Conwaylife.scala 31:34]
  wire  _T_613 = _T_612 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_614 = _T_612 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_615 = _T_612 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_616 = regs_1_3 + regs_1_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1240 = {{1'd0}, regs_1_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_617 = _T_616 + _GEN_1240; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1241 = {{2'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_618 = _T_617 + _GEN_1241; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1242 = {{3'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_619 = _T_618 + _GEN_1242; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1243 = {{4'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_620 = _T_619 + _GEN_1243; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1244 = {{5'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_621 = _T_620 + _GEN_1244; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1245 = {{6'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_622 = _T_621 + _GEN_1245; // @[Conwaylife.scala 31:34]
  wire  _T_623 = _T_622 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_624 = _T_622 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_625 = _T_622 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_626 = regs_1_4 + regs_1_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1246 = {{1'd0}, regs_1_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_627 = _T_626 + _GEN_1246; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1247 = {{2'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_628 = _T_627 + _GEN_1247; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1248 = {{3'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_629 = _T_628 + _GEN_1248; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1249 = {{4'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_630 = _T_629 + _GEN_1249; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1250 = {{5'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_631 = _T_630 + _GEN_1250; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1251 = {{6'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_632 = _T_631 + _GEN_1251; // @[Conwaylife.scala 31:34]
  wire  _T_633 = _T_632 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_634 = _T_632 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_635 = _T_632 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_636 = regs_1_5 + regs_1_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1252 = {{1'd0}, regs_1_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_637 = _T_636 + _GEN_1252; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1253 = {{2'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_638 = _T_637 + _GEN_1253; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1254 = {{3'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_639 = _T_638 + _GEN_1254; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1255 = {{4'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_640 = _T_639 + _GEN_1255; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1256 = {{5'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_641 = _T_640 + _GEN_1256; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1257 = {{6'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_642 = _T_641 + _GEN_1257; // @[Conwaylife.scala 31:34]
  wire  _T_643 = _T_642 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_644 = _T_642 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_645 = _T_642 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_646 = regs_1_6 + regs_1_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1258 = {{1'd0}, regs_1_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_647 = _T_646 + _GEN_1258; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1259 = {{2'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_648 = _T_647 + _GEN_1259; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1260 = {{3'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_649 = _T_648 + _GEN_1260; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1261 = {{4'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_650 = _T_649 + _GEN_1261; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1262 = {{5'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_651 = _T_650 + _GEN_1262; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1263 = {{6'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_652 = _T_651 + _GEN_1263; // @[Conwaylife.scala 31:34]
  wire  _T_653 = _T_652 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_654 = _T_652 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_655 = _T_652 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_656 = regs_1_7 + regs_1_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1264 = {{1'd0}, regs_1_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_657 = _T_656 + _GEN_1264; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1265 = {{2'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_658 = _T_657 + _GEN_1265; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1266 = {{3'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_659 = _T_658 + _GEN_1266; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1267 = {{4'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_660 = _T_659 + _GEN_1267; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1268 = {{5'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_661 = _T_660 + _GEN_1268; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1269 = {{6'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_662 = _T_661 + _GEN_1269; // @[Conwaylife.scala 31:34]
  wire  _T_663 = _T_662 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_664 = _T_662 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_665 = _T_662 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_666 = regs_1_8 + regs_1_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1270 = {{1'd0}, regs_1_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_667 = _T_666 + _GEN_1270; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1271 = {{2'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_668 = _T_667 + _GEN_1271; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1272 = {{3'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_669 = _T_668 + _GEN_1272; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1273 = {{4'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_670 = _T_669 + _GEN_1273; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1274 = {{5'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_671 = _T_670 + _GEN_1274; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1275 = {{6'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_672 = _T_671 + _GEN_1275; // @[Conwaylife.scala 31:34]
  wire  _T_673 = _T_672 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_674 = _T_672 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_675 = _T_672 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_676 = regs_1_9 + regs_1_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1276 = {{1'd0}, regs_1_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_677 = _T_676 + _GEN_1276; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1277 = {{2'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_678 = _T_677 + _GEN_1277; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1278 = {{3'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_679 = _T_678 + _GEN_1278; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1279 = {{4'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_680 = _T_679 + _GEN_1279; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1280 = {{5'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_681 = _T_680 + _GEN_1280; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1281 = {{6'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_682 = _T_681 + _GEN_1281; // @[Conwaylife.scala 31:34]
  wire  _T_683 = _T_682 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_684 = _T_682 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_685 = _T_682 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_686 = regs_1_10 + regs_1_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1282 = {{1'd0}, regs_1_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_687 = _T_686 + _GEN_1282; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1283 = {{2'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_688 = _T_687 + _GEN_1283; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1284 = {{3'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_689 = _T_688 + _GEN_1284; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1285 = {{4'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_690 = _T_689 + _GEN_1285; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1286 = {{5'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_691 = _T_690 + _GEN_1286; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1287 = {{6'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_692 = _T_691 + _GEN_1287; // @[Conwaylife.scala 31:34]
  wire  _T_693 = _T_692 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_694 = _T_692 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_695 = _T_692 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_696 = regs_1_11 + regs_1_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1288 = {{1'd0}, regs_1_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_697 = _T_696 + _GEN_1288; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1289 = {{2'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_698 = _T_697 + _GEN_1289; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1290 = {{3'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_699 = _T_698 + _GEN_1290; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1291 = {{4'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_700 = _T_699 + _GEN_1291; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1292 = {{5'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_701 = _T_700 + _GEN_1292; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1293 = {{6'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_702 = _T_701 + _GEN_1293; // @[Conwaylife.scala 31:34]
  wire  _T_703 = _T_702 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_704 = _T_702 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_705 = _T_702 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_706 = regs_1_12 + regs_1_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1294 = {{1'd0}, regs_1_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_707 = _T_706 + _GEN_1294; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1295 = {{2'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_708 = _T_707 + _GEN_1295; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1296 = {{3'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_709 = _T_708 + _GEN_1296; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1297 = {{4'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_710 = _T_709 + _GEN_1297; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1298 = {{5'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_711 = _T_710 + _GEN_1298; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1299 = {{6'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_712 = _T_711 + _GEN_1299; // @[Conwaylife.scala 31:34]
  wire  _T_713 = _T_712 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_714 = _T_712 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_715 = _T_712 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_716 = regs_1_13 + regs_1_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1300 = {{1'd0}, regs_1_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_717 = _T_716 + _GEN_1300; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1301 = {{2'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_718 = _T_717 + _GEN_1301; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1302 = {{3'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_719 = _T_718 + _GEN_1302; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1303 = {{4'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_720 = _T_719 + _GEN_1303; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1304 = {{5'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_721 = _T_720 + _GEN_1304; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1305 = {{6'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_722 = _T_721 + _GEN_1305; // @[Conwaylife.scala 31:34]
  wire  _T_723 = _T_722 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_724 = _T_722 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_725 = _T_722 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_726 = regs_1_14 + regs_1_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1306 = {{1'd0}, regs_1_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_727 = _T_726 + _GEN_1306; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1307 = {{2'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_728 = _T_727 + _GEN_1307; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1308 = {{3'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_729 = _T_728 + _GEN_1308; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1309 = {{4'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_730 = _T_729 + _GEN_1309; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1310 = {{5'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_731 = _T_730 + _GEN_1310; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1311 = {{6'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_732 = _T_731 + _GEN_1311; // @[Conwaylife.scala 31:34]
  wire  _T_733 = _T_732 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_734 = _T_732 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_735 = _T_732 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_736 = regs_2_15 + regs_2_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1312 = {{1'd0}, regs_2_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_737 = _T_736 + _GEN_1312; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1313 = {{2'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_738 = _T_737 + _GEN_1313; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1314 = {{3'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_739 = _T_738 + _GEN_1314; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1315 = {{4'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_740 = _T_739 + _GEN_1315; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1316 = {{5'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_741 = _T_740 + _GEN_1316; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1317 = {{6'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_742 = _T_741 + _GEN_1317; // @[Conwaylife.scala 31:34]
  wire  _T_743 = _T_742 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_744 = _T_742 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_745 = _T_742 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_746 = regs_2_0 + regs_2_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1318 = {{1'd0}, regs_2_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_747 = _T_746 + _GEN_1318; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1319 = {{2'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_748 = _T_747 + _GEN_1319; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1320 = {{3'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_749 = _T_748 + _GEN_1320; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1321 = {{4'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_750 = _T_749 + _GEN_1321; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1322 = {{5'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_751 = _T_750 + _GEN_1322; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1323 = {{6'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_752 = _T_751 + _GEN_1323; // @[Conwaylife.scala 31:34]
  wire  _T_753 = _T_752 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_754 = _T_752 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_755 = _T_752 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_756 = regs_2_1 + regs_2_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1324 = {{1'd0}, regs_2_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_757 = _T_756 + _GEN_1324; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1325 = {{2'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_758 = _T_757 + _GEN_1325; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1326 = {{3'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_759 = _T_758 + _GEN_1326; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1327 = {{4'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_760 = _T_759 + _GEN_1327; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1328 = {{5'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_761 = _T_760 + _GEN_1328; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1329 = {{6'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_762 = _T_761 + _GEN_1329; // @[Conwaylife.scala 31:34]
  wire  _T_763 = _T_762 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_764 = _T_762 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_765 = _T_762 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_766 = regs_2_2 + regs_2_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1330 = {{1'd0}, regs_2_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_767 = _T_766 + _GEN_1330; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1331 = {{2'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_768 = _T_767 + _GEN_1331; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1332 = {{3'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_769 = _T_768 + _GEN_1332; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1333 = {{4'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_770 = _T_769 + _GEN_1333; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1334 = {{5'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_771 = _T_770 + _GEN_1334; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1335 = {{6'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_772 = _T_771 + _GEN_1335; // @[Conwaylife.scala 31:34]
  wire  _T_773 = _T_772 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_774 = _T_772 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_775 = _T_772 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_776 = regs_2_3 + regs_2_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1336 = {{1'd0}, regs_2_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_777 = _T_776 + _GEN_1336; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1337 = {{2'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_778 = _T_777 + _GEN_1337; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1338 = {{3'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_779 = _T_778 + _GEN_1338; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1339 = {{4'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_780 = _T_779 + _GEN_1339; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1340 = {{5'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_781 = _T_780 + _GEN_1340; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1341 = {{6'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_782 = _T_781 + _GEN_1341; // @[Conwaylife.scala 31:34]
  wire  _T_783 = _T_782 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_784 = _T_782 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_785 = _T_782 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_786 = regs_2_4 + regs_2_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1342 = {{1'd0}, regs_2_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_787 = _T_786 + _GEN_1342; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1343 = {{2'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_788 = _T_787 + _GEN_1343; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1344 = {{3'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_789 = _T_788 + _GEN_1344; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1345 = {{4'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_790 = _T_789 + _GEN_1345; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1346 = {{5'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_791 = _T_790 + _GEN_1346; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1347 = {{6'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_792 = _T_791 + _GEN_1347; // @[Conwaylife.scala 31:34]
  wire  _T_793 = _T_792 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_794 = _T_792 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_795 = _T_792 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_796 = regs_2_5 + regs_2_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1348 = {{1'd0}, regs_2_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_797 = _T_796 + _GEN_1348; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1349 = {{2'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_798 = _T_797 + _GEN_1349; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1350 = {{3'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_799 = _T_798 + _GEN_1350; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1351 = {{4'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_800 = _T_799 + _GEN_1351; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1352 = {{5'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_801 = _T_800 + _GEN_1352; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1353 = {{6'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_802 = _T_801 + _GEN_1353; // @[Conwaylife.scala 31:34]
  wire  _T_803 = _T_802 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_804 = _T_802 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_805 = _T_802 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_806 = regs_2_6 + regs_2_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1354 = {{1'd0}, regs_2_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_807 = _T_806 + _GEN_1354; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1355 = {{2'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_808 = _T_807 + _GEN_1355; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1356 = {{3'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_809 = _T_808 + _GEN_1356; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1357 = {{4'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_810 = _T_809 + _GEN_1357; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1358 = {{5'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_811 = _T_810 + _GEN_1358; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1359 = {{6'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_812 = _T_811 + _GEN_1359; // @[Conwaylife.scala 31:34]
  wire  _T_813 = _T_812 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_814 = _T_812 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_815 = _T_812 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_816 = regs_2_7 + regs_2_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1360 = {{1'd0}, regs_2_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_817 = _T_816 + _GEN_1360; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1361 = {{2'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_818 = _T_817 + _GEN_1361; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1362 = {{3'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_819 = _T_818 + _GEN_1362; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1363 = {{4'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_820 = _T_819 + _GEN_1363; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1364 = {{5'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_821 = _T_820 + _GEN_1364; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1365 = {{6'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_822 = _T_821 + _GEN_1365; // @[Conwaylife.scala 31:34]
  wire  _T_823 = _T_822 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_824 = _T_822 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_825 = _T_822 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_826 = regs_2_8 + regs_2_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1366 = {{1'd0}, regs_2_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_827 = _T_826 + _GEN_1366; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1367 = {{2'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_828 = _T_827 + _GEN_1367; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1368 = {{3'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_829 = _T_828 + _GEN_1368; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1369 = {{4'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_830 = _T_829 + _GEN_1369; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1370 = {{5'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_831 = _T_830 + _GEN_1370; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1371 = {{6'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_832 = _T_831 + _GEN_1371; // @[Conwaylife.scala 31:34]
  wire  _T_833 = _T_832 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_834 = _T_832 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_835 = _T_832 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_836 = regs_2_9 + regs_2_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1372 = {{1'd0}, regs_2_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_837 = _T_836 + _GEN_1372; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1373 = {{2'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_838 = _T_837 + _GEN_1373; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1374 = {{3'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_839 = _T_838 + _GEN_1374; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1375 = {{4'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_840 = _T_839 + _GEN_1375; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1376 = {{5'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_841 = _T_840 + _GEN_1376; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1377 = {{6'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_842 = _T_841 + _GEN_1377; // @[Conwaylife.scala 31:34]
  wire  _T_843 = _T_842 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_844 = _T_842 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_845 = _T_842 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_846 = regs_2_10 + regs_2_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1378 = {{1'd0}, regs_2_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_847 = _T_846 + _GEN_1378; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1379 = {{2'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_848 = _T_847 + _GEN_1379; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1380 = {{3'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_849 = _T_848 + _GEN_1380; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1381 = {{4'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_850 = _T_849 + _GEN_1381; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1382 = {{5'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_851 = _T_850 + _GEN_1382; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1383 = {{6'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_852 = _T_851 + _GEN_1383; // @[Conwaylife.scala 31:34]
  wire  _T_853 = _T_852 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_854 = _T_852 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_855 = _T_852 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_856 = regs_2_11 + regs_2_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1384 = {{1'd0}, regs_2_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_857 = _T_856 + _GEN_1384; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1385 = {{2'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_858 = _T_857 + _GEN_1385; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1386 = {{3'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_859 = _T_858 + _GEN_1386; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1387 = {{4'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_860 = _T_859 + _GEN_1387; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1388 = {{5'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_861 = _T_860 + _GEN_1388; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1389 = {{6'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_862 = _T_861 + _GEN_1389; // @[Conwaylife.scala 31:34]
  wire  _T_863 = _T_862 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_864 = _T_862 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_865 = _T_862 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_866 = regs_2_12 + regs_2_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1390 = {{1'd0}, regs_2_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_867 = _T_866 + _GEN_1390; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1391 = {{2'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_868 = _T_867 + _GEN_1391; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1392 = {{3'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_869 = _T_868 + _GEN_1392; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1393 = {{4'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_870 = _T_869 + _GEN_1393; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1394 = {{5'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_871 = _T_870 + _GEN_1394; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1395 = {{6'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_872 = _T_871 + _GEN_1395; // @[Conwaylife.scala 31:34]
  wire  _T_873 = _T_872 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_874 = _T_872 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_875 = _T_872 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_876 = regs_2_13 + regs_2_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1396 = {{1'd0}, regs_2_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_877 = _T_876 + _GEN_1396; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1397 = {{2'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_878 = _T_877 + _GEN_1397; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1398 = {{3'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_879 = _T_878 + _GEN_1398; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1399 = {{4'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_880 = _T_879 + _GEN_1399; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1400 = {{5'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_881 = _T_880 + _GEN_1400; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1401 = {{6'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_882 = _T_881 + _GEN_1401; // @[Conwaylife.scala 31:34]
  wire  _T_883 = _T_882 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_884 = _T_882 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_885 = _T_882 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_886 = regs_2_14 + regs_2_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1402 = {{1'd0}, regs_2_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_887 = _T_886 + _GEN_1402; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1403 = {{2'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_888 = _T_887 + _GEN_1403; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1404 = {{3'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_889 = _T_888 + _GEN_1404; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1405 = {{4'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_890 = _T_889 + _GEN_1405; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1406 = {{5'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_891 = _T_890 + _GEN_1406; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1407 = {{6'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_892 = _T_891 + _GEN_1407; // @[Conwaylife.scala 31:34]
  wire  _T_893 = _T_892 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_894 = _T_892 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_895 = _T_892 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_896 = regs_3_15 + regs_3_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1408 = {{1'd0}, regs_3_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_897 = _T_896 + _GEN_1408; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1409 = {{2'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_898 = _T_897 + _GEN_1409; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1410 = {{3'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_899 = _T_898 + _GEN_1410; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1411 = {{4'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_900 = _T_899 + _GEN_1411; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1412 = {{5'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_901 = _T_900 + _GEN_1412; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1413 = {{6'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_902 = _T_901 + _GEN_1413; // @[Conwaylife.scala 31:34]
  wire  _T_903 = _T_902 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_904 = _T_902 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_905 = _T_902 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_906 = regs_3_0 + regs_3_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1414 = {{1'd0}, regs_3_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_907 = _T_906 + _GEN_1414; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1415 = {{2'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_908 = _T_907 + _GEN_1415; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1416 = {{3'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_909 = _T_908 + _GEN_1416; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1417 = {{4'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_910 = _T_909 + _GEN_1417; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1418 = {{5'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_911 = _T_910 + _GEN_1418; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1419 = {{6'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_912 = _T_911 + _GEN_1419; // @[Conwaylife.scala 31:34]
  wire  _T_913 = _T_912 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_914 = _T_912 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_915 = _T_912 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_916 = regs_3_1 + regs_3_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1420 = {{1'd0}, regs_3_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_917 = _T_916 + _GEN_1420; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1421 = {{2'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_918 = _T_917 + _GEN_1421; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1422 = {{3'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_919 = _T_918 + _GEN_1422; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1423 = {{4'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_920 = _T_919 + _GEN_1423; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1424 = {{5'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_921 = _T_920 + _GEN_1424; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1425 = {{6'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_922 = _T_921 + _GEN_1425; // @[Conwaylife.scala 31:34]
  wire  _T_923 = _T_922 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_924 = _T_922 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_925 = _T_922 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_926 = regs_3_2 + regs_3_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1426 = {{1'd0}, regs_3_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_927 = _T_926 + _GEN_1426; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1427 = {{2'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_928 = _T_927 + _GEN_1427; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1428 = {{3'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_929 = _T_928 + _GEN_1428; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1429 = {{4'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_930 = _T_929 + _GEN_1429; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1430 = {{5'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_931 = _T_930 + _GEN_1430; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1431 = {{6'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_932 = _T_931 + _GEN_1431; // @[Conwaylife.scala 31:34]
  wire  _T_933 = _T_932 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_934 = _T_932 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_935 = _T_932 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_936 = regs_3_3 + regs_3_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1432 = {{1'd0}, regs_3_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_937 = _T_936 + _GEN_1432; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1433 = {{2'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_938 = _T_937 + _GEN_1433; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1434 = {{3'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_939 = _T_938 + _GEN_1434; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1435 = {{4'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_940 = _T_939 + _GEN_1435; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1436 = {{5'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_941 = _T_940 + _GEN_1436; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1437 = {{6'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_942 = _T_941 + _GEN_1437; // @[Conwaylife.scala 31:34]
  wire  _T_943 = _T_942 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_944 = _T_942 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_945 = _T_942 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_946 = regs_3_4 + regs_3_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1438 = {{1'd0}, regs_3_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_947 = _T_946 + _GEN_1438; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1439 = {{2'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_948 = _T_947 + _GEN_1439; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1440 = {{3'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_949 = _T_948 + _GEN_1440; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1441 = {{4'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_950 = _T_949 + _GEN_1441; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1442 = {{5'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_951 = _T_950 + _GEN_1442; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1443 = {{6'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_952 = _T_951 + _GEN_1443; // @[Conwaylife.scala 31:34]
  wire  _T_953 = _T_952 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_954 = _T_952 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_955 = _T_952 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_956 = regs_3_5 + regs_3_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1444 = {{1'd0}, regs_3_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_957 = _T_956 + _GEN_1444; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1445 = {{2'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_958 = _T_957 + _GEN_1445; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1446 = {{3'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_959 = _T_958 + _GEN_1446; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1447 = {{4'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_960 = _T_959 + _GEN_1447; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1448 = {{5'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_961 = _T_960 + _GEN_1448; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1449 = {{6'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_962 = _T_961 + _GEN_1449; // @[Conwaylife.scala 31:34]
  wire  _T_963 = _T_962 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_964 = _T_962 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_965 = _T_962 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_966 = regs_3_6 + regs_3_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1450 = {{1'd0}, regs_3_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_967 = _T_966 + _GEN_1450; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1451 = {{2'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_968 = _T_967 + _GEN_1451; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1452 = {{3'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_969 = _T_968 + _GEN_1452; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1453 = {{4'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_970 = _T_969 + _GEN_1453; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1454 = {{5'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_971 = _T_970 + _GEN_1454; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1455 = {{6'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_972 = _T_971 + _GEN_1455; // @[Conwaylife.scala 31:34]
  wire  _T_973 = _T_972 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_974 = _T_972 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_975 = _T_972 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_976 = regs_3_7 + regs_3_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1456 = {{1'd0}, regs_3_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_977 = _T_976 + _GEN_1456; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1457 = {{2'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_978 = _T_977 + _GEN_1457; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1458 = {{3'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_979 = _T_978 + _GEN_1458; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1459 = {{4'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_980 = _T_979 + _GEN_1459; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1460 = {{5'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_981 = _T_980 + _GEN_1460; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1461 = {{6'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_982 = _T_981 + _GEN_1461; // @[Conwaylife.scala 31:34]
  wire  _T_983 = _T_982 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_984 = _T_982 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_985 = _T_982 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_986 = regs_3_8 + regs_3_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1462 = {{1'd0}, regs_3_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_987 = _T_986 + _GEN_1462; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1463 = {{2'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_988 = _T_987 + _GEN_1463; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1464 = {{3'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_989 = _T_988 + _GEN_1464; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1465 = {{4'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_990 = _T_989 + _GEN_1465; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1466 = {{5'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_991 = _T_990 + _GEN_1466; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1467 = {{6'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_992 = _T_991 + _GEN_1467; // @[Conwaylife.scala 31:34]
  wire  _T_993 = _T_992 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_994 = _T_992 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_995 = _T_992 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_996 = regs_3_9 + regs_3_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1468 = {{1'd0}, regs_3_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_997 = _T_996 + _GEN_1468; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1469 = {{2'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_998 = _T_997 + _GEN_1469; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1470 = {{3'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_999 = _T_998 + _GEN_1470; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1471 = {{4'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1000 = _T_999 + _GEN_1471; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1472 = {{5'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1001 = _T_1000 + _GEN_1472; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1473 = {{6'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1002 = _T_1001 + _GEN_1473; // @[Conwaylife.scala 31:34]
  wire  _T_1003 = _T_1002 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1004 = _T_1002 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1005 = _T_1002 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1006 = regs_3_10 + regs_3_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1474 = {{1'd0}, regs_3_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1007 = _T_1006 + _GEN_1474; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1475 = {{2'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1008 = _T_1007 + _GEN_1475; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1476 = {{3'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1009 = _T_1008 + _GEN_1476; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1477 = {{4'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1010 = _T_1009 + _GEN_1477; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1478 = {{5'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1011 = _T_1010 + _GEN_1478; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1479 = {{6'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1012 = _T_1011 + _GEN_1479; // @[Conwaylife.scala 31:34]
  wire  _T_1013 = _T_1012 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1014 = _T_1012 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1015 = _T_1012 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1016 = regs_3_11 + regs_3_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1480 = {{1'd0}, regs_3_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1017 = _T_1016 + _GEN_1480; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1481 = {{2'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1018 = _T_1017 + _GEN_1481; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1482 = {{3'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1019 = _T_1018 + _GEN_1482; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1483 = {{4'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1020 = _T_1019 + _GEN_1483; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1484 = {{5'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1021 = _T_1020 + _GEN_1484; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1485 = {{6'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1022 = _T_1021 + _GEN_1485; // @[Conwaylife.scala 31:34]
  wire  _T_1023 = _T_1022 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1024 = _T_1022 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1025 = _T_1022 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1026 = regs_3_12 + regs_3_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1486 = {{1'd0}, regs_3_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1027 = _T_1026 + _GEN_1486; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1487 = {{2'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1028 = _T_1027 + _GEN_1487; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1488 = {{3'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1029 = _T_1028 + _GEN_1488; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1489 = {{4'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1030 = _T_1029 + _GEN_1489; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1490 = {{5'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1031 = _T_1030 + _GEN_1490; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1491 = {{6'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1032 = _T_1031 + _GEN_1491; // @[Conwaylife.scala 31:34]
  wire  _T_1033 = _T_1032 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1034 = _T_1032 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1035 = _T_1032 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1036 = regs_3_13 + regs_3_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1492 = {{1'd0}, regs_3_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1037 = _T_1036 + _GEN_1492; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1493 = {{2'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1038 = _T_1037 + _GEN_1493; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1494 = {{3'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1039 = _T_1038 + _GEN_1494; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1495 = {{4'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1040 = _T_1039 + _GEN_1495; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1496 = {{5'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1041 = _T_1040 + _GEN_1496; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1497 = {{6'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1042 = _T_1041 + _GEN_1497; // @[Conwaylife.scala 31:34]
  wire  _T_1043 = _T_1042 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1044 = _T_1042 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1045 = _T_1042 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1046 = regs_3_14 + regs_3_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1498 = {{1'd0}, regs_3_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1047 = _T_1046 + _GEN_1498; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1499 = {{2'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1048 = _T_1047 + _GEN_1499; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1500 = {{3'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1049 = _T_1048 + _GEN_1500; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1501 = {{4'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1050 = _T_1049 + _GEN_1501; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1502 = {{5'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1051 = _T_1050 + _GEN_1502; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1503 = {{6'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1052 = _T_1051 + _GEN_1503; // @[Conwaylife.scala 31:34]
  wire  _T_1053 = _T_1052 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1054 = _T_1052 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1055 = _T_1052 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1056 = regs_4_15 + regs_4_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1504 = {{1'd0}, regs_4_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1057 = _T_1056 + _GEN_1504; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1505 = {{2'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1058 = _T_1057 + _GEN_1505; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1506 = {{3'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1059 = _T_1058 + _GEN_1506; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1507 = {{4'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1060 = _T_1059 + _GEN_1507; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1508 = {{5'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1061 = _T_1060 + _GEN_1508; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1509 = {{6'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1062 = _T_1061 + _GEN_1509; // @[Conwaylife.scala 31:34]
  wire  _T_1063 = _T_1062 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1064 = _T_1062 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1065 = _T_1062 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1066 = regs_4_0 + regs_4_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1510 = {{1'd0}, regs_4_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1067 = _T_1066 + _GEN_1510; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1511 = {{2'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1068 = _T_1067 + _GEN_1511; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1512 = {{3'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1069 = _T_1068 + _GEN_1512; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1513 = {{4'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1070 = _T_1069 + _GEN_1513; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1514 = {{5'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1071 = _T_1070 + _GEN_1514; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1515 = {{6'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1072 = _T_1071 + _GEN_1515; // @[Conwaylife.scala 31:34]
  wire  _T_1073 = _T_1072 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1074 = _T_1072 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1075 = _T_1072 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1076 = regs_4_1 + regs_4_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1516 = {{1'd0}, regs_4_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1077 = _T_1076 + _GEN_1516; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1517 = {{2'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1078 = _T_1077 + _GEN_1517; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1518 = {{3'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1079 = _T_1078 + _GEN_1518; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1519 = {{4'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1080 = _T_1079 + _GEN_1519; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1520 = {{5'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1081 = _T_1080 + _GEN_1520; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1521 = {{6'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1082 = _T_1081 + _GEN_1521; // @[Conwaylife.scala 31:34]
  wire  _T_1083 = _T_1082 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1084 = _T_1082 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1085 = _T_1082 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1086 = regs_4_2 + regs_4_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1522 = {{1'd0}, regs_4_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1087 = _T_1086 + _GEN_1522; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1523 = {{2'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1088 = _T_1087 + _GEN_1523; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1524 = {{3'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1089 = _T_1088 + _GEN_1524; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1525 = {{4'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1090 = _T_1089 + _GEN_1525; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1526 = {{5'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1091 = _T_1090 + _GEN_1526; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1527 = {{6'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1092 = _T_1091 + _GEN_1527; // @[Conwaylife.scala 31:34]
  wire  _T_1093 = _T_1092 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1094 = _T_1092 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1095 = _T_1092 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1096 = regs_4_3 + regs_4_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1528 = {{1'd0}, regs_4_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1097 = _T_1096 + _GEN_1528; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1529 = {{2'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1098 = _T_1097 + _GEN_1529; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1530 = {{3'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1099 = _T_1098 + _GEN_1530; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1531 = {{4'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1100 = _T_1099 + _GEN_1531; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1532 = {{5'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1101 = _T_1100 + _GEN_1532; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1533 = {{6'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1102 = _T_1101 + _GEN_1533; // @[Conwaylife.scala 31:34]
  wire  _T_1103 = _T_1102 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1104 = _T_1102 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1105 = _T_1102 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1106 = regs_4_4 + regs_4_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1534 = {{1'd0}, regs_4_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1107 = _T_1106 + _GEN_1534; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1535 = {{2'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1108 = _T_1107 + _GEN_1535; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1536 = {{3'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1109 = _T_1108 + _GEN_1536; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1537 = {{4'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1110 = _T_1109 + _GEN_1537; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1538 = {{5'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1111 = _T_1110 + _GEN_1538; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1539 = {{6'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1112 = _T_1111 + _GEN_1539; // @[Conwaylife.scala 31:34]
  wire  _T_1113 = _T_1112 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1114 = _T_1112 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1115 = _T_1112 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1116 = regs_4_5 + regs_4_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1540 = {{1'd0}, regs_4_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1117 = _T_1116 + _GEN_1540; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1541 = {{2'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1118 = _T_1117 + _GEN_1541; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1542 = {{3'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1119 = _T_1118 + _GEN_1542; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1543 = {{4'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1120 = _T_1119 + _GEN_1543; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1544 = {{5'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1121 = _T_1120 + _GEN_1544; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1545 = {{6'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1122 = _T_1121 + _GEN_1545; // @[Conwaylife.scala 31:34]
  wire  _T_1123 = _T_1122 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1124 = _T_1122 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1125 = _T_1122 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1126 = regs_4_6 + regs_4_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1546 = {{1'd0}, regs_4_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1127 = _T_1126 + _GEN_1546; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1547 = {{2'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1128 = _T_1127 + _GEN_1547; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1548 = {{3'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1129 = _T_1128 + _GEN_1548; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1549 = {{4'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1130 = _T_1129 + _GEN_1549; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1550 = {{5'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1131 = _T_1130 + _GEN_1550; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1551 = {{6'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1132 = _T_1131 + _GEN_1551; // @[Conwaylife.scala 31:34]
  wire  _T_1133 = _T_1132 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1134 = _T_1132 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1135 = _T_1132 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1136 = regs_4_7 + regs_4_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1552 = {{1'd0}, regs_4_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1137 = _T_1136 + _GEN_1552; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1553 = {{2'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1138 = _T_1137 + _GEN_1553; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1554 = {{3'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1139 = _T_1138 + _GEN_1554; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1555 = {{4'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1140 = _T_1139 + _GEN_1555; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1556 = {{5'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1141 = _T_1140 + _GEN_1556; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1557 = {{6'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1142 = _T_1141 + _GEN_1557; // @[Conwaylife.scala 31:34]
  wire  _T_1143 = _T_1142 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1144 = _T_1142 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1145 = _T_1142 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1146 = regs_4_8 + regs_4_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1558 = {{1'd0}, regs_4_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1147 = _T_1146 + _GEN_1558; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1559 = {{2'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1148 = _T_1147 + _GEN_1559; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1560 = {{3'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1149 = _T_1148 + _GEN_1560; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1561 = {{4'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1150 = _T_1149 + _GEN_1561; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1562 = {{5'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1151 = _T_1150 + _GEN_1562; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1563 = {{6'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1152 = _T_1151 + _GEN_1563; // @[Conwaylife.scala 31:34]
  wire  _T_1153 = _T_1152 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1154 = _T_1152 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1155 = _T_1152 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1156 = regs_4_9 + regs_4_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1564 = {{1'd0}, regs_4_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1157 = _T_1156 + _GEN_1564; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1565 = {{2'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1158 = _T_1157 + _GEN_1565; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1566 = {{3'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1159 = _T_1158 + _GEN_1566; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1567 = {{4'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1160 = _T_1159 + _GEN_1567; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1568 = {{5'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1161 = _T_1160 + _GEN_1568; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1569 = {{6'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1162 = _T_1161 + _GEN_1569; // @[Conwaylife.scala 31:34]
  wire  _T_1163 = _T_1162 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1164 = _T_1162 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1165 = _T_1162 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1166 = regs_4_10 + regs_4_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1570 = {{1'd0}, regs_4_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1167 = _T_1166 + _GEN_1570; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1571 = {{2'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1168 = _T_1167 + _GEN_1571; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1572 = {{3'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1169 = _T_1168 + _GEN_1572; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1573 = {{4'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1170 = _T_1169 + _GEN_1573; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1574 = {{5'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1171 = _T_1170 + _GEN_1574; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1575 = {{6'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1172 = _T_1171 + _GEN_1575; // @[Conwaylife.scala 31:34]
  wire  _T_1173 = _T_1172 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1174 = _T_1172 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1175 = _T_1172 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1176 = regs_4_11 + regs_4_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1576 = {{1'd0}, regs_4_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1177 = _T_1176 + _GEN_1576; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1577 = {{2'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1178 = _T_1177 + _GEN_1577; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1578 = {{3'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1179 = _T_1178 + _GEN_1578; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1579 = {{4'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1180 = _T_1179 + _GEN_1579; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1580 = {{5'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1181 = _T_1180 + _GEN_1580; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1581 = {{6'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1182 = _T_1181 + _GEN_1581; // @[Conwaylife.scala 31:34]
  wire  _T_1183 = _T_1182 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1184 = _T_1182 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1185 = _T_1182 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1186 = regs_4_12 + regs_4_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1582 = {{1'd0}, regs_4_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1187 = _T_1186 + _GEN_1582; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1583 = {{2'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1188 = _T_1187 + _GEN_1583; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1584 = {{3'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1189 = _T_1188 + _GEN_1584; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1585 = {{4'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1190 = _T_1189 + _GEN_1585; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1586 = {{5'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1191 = _T_1190 + _GEN_1586; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1587 = {{6'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1192 = _T_1191 + _GEN_1587; // @[Conwaylife.scala 31:34]
  wire  _T_1193 = _T_1192 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1194 = _T_1192 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1195 = _T_1192 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1196 = regs_4_13 + regs_4_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1588 = {{1'd0}, regs_4_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1197 = _T_1196 + _GEN_1588; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1589 = {{2'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1198 = _T_1197 + _GEN_1589; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1590 = {{3'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1199 = _T_1198 + _GEN_1590; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1591 = {{4'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1200 = _T_1199 + _GEN_1591; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1592 = {{5'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1201 = _T_1200 + _GEN_1592; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1593 = {{6'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1202 = _T_1201 + _GEN_1593; // @[Conwaylife.scala 31:34]
  wire  _T_1203 = _T_1202 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1204 = _T_1202 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1205 = _T_1202 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1206 = regs_4_14 + regs_4_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1594 = {{1'd0}, regs_4_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1207 = _T_1206 + _GEN_1594; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1595 = {{2'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1208 = _T_1207 + _GEN_1595; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1596 = {{3'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1209 = _T_1208 + _GEN_1596; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1597 = {{4'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1210 = _T_1209 + _GEN_1597; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1598 = {{5'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1211 = _T_1210 + _GEN_1598; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1599 = {{6'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1212 = _T_1211 + _GEN_1599; // @[Conwaylife.scala 31:34]
  wire  _T_1213 = _T_1212 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1214 = _T_1212 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1215 = _T_1212 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1216 = regs_5_15 + regs_5_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1600 = {{1'd0}, regs_5_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1217 = _T_1216 + _GEN_1600; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1601 = {{2'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1218 = _T_1217 + _GEN_1601; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1602 = {{3'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1219 = _T_1218 + _GEN_1602; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1603 = {{4'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1220 = _T_1219 + _GEN_1603; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1604 = {{5'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1221 = _T_1220 + _GEN_1604; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1605 = {{6'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1222 = _T_1221 + _GEN_1605; // @[Conwaylife.scala 31:34]
  wire  _T_1223 = _T_1222 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1224 = _T_1222 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1225 = _T_1222 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1226 = regs_5_0 + regs_5_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1606 = {{1'd0}, regs_5_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1227 = _T_1226 + _GEN_1606; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1607 = {{2'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1228 = _T_1227 + _GEN_1607; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1608 = {{3'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1229 = _T_1228 + _GEN_1608; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1609 = {{4'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1230 = _T_1229 + _GEN_1609; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1610 = {{5'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1231 = _T_1230 + _GEN_1610; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1611 = {{6'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1232 = _T_1231 + _GEN_1611; // @[Conwaylife.scala 31:34]
  wire  _T_1233 = _T_1232 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1234 = _T_1232 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1235 = _T_1232 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1236 = regs_5_1 + regs_5_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1612 = {{1'd0}, regs_5_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1237 = _T_1236 + _GEN_1612; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1613 = {{2'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1238 = _T_1237 + _GEN_1613; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1614 = {{3'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1239 = _T_1238 + _GEN_1614; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1615 = {{4'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1240 = _T_1239 + _GEN_1615; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1616 = {{5'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1241 = _T_1240 + _GEN_1616; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1617 = {{6'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1242 = _T_1241 + _GEN_1617; // @[Conwaylife.scala 31:34]
  wire  _T_1243 = _T_1242 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1244 = _T_1242 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1245 = _T_1242 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1246 = regs_5_2 + regs_5_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1618 = {{1'd0}, regs_5_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1247 = _T_1246 + _GEN_1618; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1619 = {{2'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1248 = _T_1247 + _GEN_1619; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1620 = {{3'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1249 = _T_1248 + _GEN_1620; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1621 = {{4'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1250 = _T_1249 + _GEN_1621; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1622 = {{5'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1251 = _T_1250 + _GEN_1622; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1623 = {{6'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1252 = _T_1251 + _GEN_1623; // @[Conwaylife.scala 31:34]
  wire  _T_1253 = _T_1252 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1254 = _T_1252 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1255 = _T_1252 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1256 = regs_5_3 + regs_5_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1624 = {{1'd0}, regs_5_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1257 = _T_1256 + _GEN_1624; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1625 = {{2'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1258 = _T_1257 + _GEN_1625; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1626 = {{3'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1259 = _T_1258 + _GEN_1626; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1627 = {{4'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1260 = _T_1259 + _GEN_1627; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1628 = {{5'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1261 = _T_1260 + _GEN_1628; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1629 = {{6'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1262 = _T_1261 + _GEN_1629; // @[Conwaylife.scala 31:34]
  wire  _T_1263 = _T_1262 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1264 = _T_1262 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1265 = _T_1262 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1266 = regs_5_4 + regs_5_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1630 = {{1'd0}, regs_5_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1267 = _T_1266 + _GEN_1630; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1631 = {{2'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1268 = _T_1267 + _GEN_1631; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1632 = {{3'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1269 = _T_1268 + _GEN_1632; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1633 = {{4'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1270 = _T_1269 + _GEN_1633; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1634 = {{5'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1271 = _T_1270 + _GEN_1634; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1635 = {{6'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1272 = _T_1271 + _GEN_1635; // @[Conwaylife.scala 31:34]
  wire  _T_1273 = _T_1272 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1274 = _T_1272 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1275 = _T_1272 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1276 = regs_5_5 + regs_5_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1636 = {{1'd0}, regs_5_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1277 = _T_1276 + _GEN_1636; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1637 = {{2'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1278 = _T_1277 + _GEN_1637; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1638 = {{3'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1279 = _T_1278 + _GEN_1638; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1639 = {{4'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1280 = _T_1279 + _GEN_1639; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1640 = {{5'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1281 = _T_1280 + _GEN_1640; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1641 = {{6'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1282 = _T_1281 + _GEN_1641; // @[Conwaylife.scala 31:34]
  wire  _T_1283 = _T_1282 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1284 = _T_1282 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1285 = _T_1282 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1286 = regs_5_6 + regs_5_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1642 = {{1'd0}, regs_5_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1287 = _T_1286 + _GEN_1642; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1643 = {{2'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1288 = _T_1287 + _GEN_1643; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1644 = {{3'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1289 = _T_1288 + _GEN_1644; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1645 = {{4'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1290 = _T_1289 + _GEN_1645; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1646 = {{5'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1291 = _T_1290 + _GEN_1646; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1647 = {{6'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1292 = _T_1291 + _GEN_1647; // @[Conwaylife.scala 31:34]
  wire  _T_1293 = _T_1292 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1294 = _T_1292 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1295 = _T_1292 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1296 = regs_5_7 + regs_5_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1648 = {{1'd0}, regs_5_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1297 = _T_1296 + _GEN_1648; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1649 = {{2'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1298 = _T_1297 + _GEN_1649; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1650 = {{3'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1299 = _T_1298 + _GEN_1650; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1651 = {{4'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1300 = _T_1299 + _GEN_1651; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1652 = {{5'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1301 = _T_1300 + _GEN_1652; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1653 = {{6'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1302 = _T_1301 + _GEN_1653; // @[Conwaylife.scala 31:34]
  wire  _T_1303 = _T_1302 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1304 = _T_1302 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1305 = _T_1302 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1306 = regs_5_8 + regs_5_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1654 = {{1'd0}, regs_5_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1307 = _T_1306 + _GEN_1654; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1655 = {{2'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1308 = _T_1307 + _GEN_1655; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1656 = {{3'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1309 = _T_1308 + _GEN_1656; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1657 = {{4'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1310 = _T_1309 + _GEN_1657; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1658 = {{5'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1311 = _T_1310 + _GEN_1658; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1659 = {{6'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1312 = _T_1311 + _GEN_1659; // @[Conwaylife.scala 31:34]
  wire  _T_1313 = _T_1312 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1314 = _T_1312 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1315 = _T_1312 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1316 = regs_5_9 + regs_5_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1660 = {{1'd0}, regs_5_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1317 = _T_1316 + _GEN_1660; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1661 = {{2'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1318 = _T_1317 + _GEN_1661; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1662 = {{3'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1319 = _T_1318 + _GEN_1662; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1663 = {{4'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1320 = _T_1319 + _GEN_1663; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1664 = {{5'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1321 = _T_1320 + _GEN_1664; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1665 = {{6'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1322 = _T_1321 + _GEN_1665; // @[Conwaylife.scala 31:34]
  wire  _T_1323 = _T_1322 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1324 = _T_1322 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1325 = _T_1322 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1326 = regs_5_10 + regs_5_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1666 = {{1'd0}, regs_5_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1327 = _T_1326 + _GEN_1666; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1667 = {{2'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1328 = _T_1327 + _GEN_1667; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1668 = {{3'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1329 = _T_1328 + _GEN_1668; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1669 = {{4'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1330 = _T_1329 + _GEN_1669; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1670 = {{5'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1331 = _T_1330 + _GEN_1670; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1671 = {{6'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1332 = _T_1331 + _GEN_1671; // @[Conwaylife.scala 31:34]
  wire  _T_1333 = _T_1332 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1334 = _T_1332 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1335 = _T_1332 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1336 = regs_5_11 + regs_5_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1672 = {{1'd0}, regs_5_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1337 = _T_1336 + _GEN_1672; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1673 = {{2'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1338 = _T_1337 + _GEN_1673; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1674 = {{3'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1339 = _T_1338 + _GEN_1674; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1675 = {{4'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1340 = _T_1339 + _GEN_1675; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1676 = {{5'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1341 = _T_1340 + _GEN_1676; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1677 = {{6'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1342 = _T_1341 + _GEN_1677; // @[Conwaylife.scala 31:34]
  wire  _T_1343 = _T_1342 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1344 = _T_1342 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1345 = _T_1342 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1346 = regs_5_12 + regs_5_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1678 = {{1'd0}, regs_5_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1347 = _T_1346 + _GEN_1678; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1679 = {{2'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1348 = _T_1347 + _GEN_1679; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1680 = {{3'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1349 = _T_1348 + _GEN_1680; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1681 = {{4'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1350 = _T_1349 + _GEN_1681; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1682 = {{5'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1351 = _T_1350 + _GEN_1682; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1683 = {{6'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1352 = _T_1351 + _GEN_1683; // @[Conwaylife.scala 31:34]
  wire  _T_1353 = _T_1352 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1354 = _T_1352 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1355 = _T_1352 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1356 = regs_5_13 + regs_5_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1684 = {{1'd0}, regs_5_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1357 = _T_1356 + _GEN_1684; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1685 = {{2'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1358 = _T_1357 + _GEN_1685; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1686 = {{3'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1359 = _T_1358 + _GEN_1686; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1687 = {{4'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1360 = _T_1359 + _GEN_1687; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1688 = {{5'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1361 = _T_1360 + _GEN_1688; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1689 = {{6'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1362 = _T_1361 + _GEN_1689; // @[Conwaylife.scala 31:34]
  wire  _T_1363 = _T_1362 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1364 = _T_1362 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1365 = _T_1362 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1366 = regs_5_14 + regs_5_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1690 = {{1'd0}, regs_5_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1367 = _T_1366 + _GEN_1690; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1691 = {{2'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1368 = _T_1367 + _GEN_1691; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1692 = {{3'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1369 = _T_1368 + _GEN_1692; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1693 = {{4'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1370 = _T_1369 + _GEN_1693; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1694 = {{5'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1371 = _T_1370 + _GEN_1694; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1695 = {{6'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1372 = _T_1371 + _GEN_1695; // @[Conwaylife.scala 31:34]
  wire  _T_1373 = _T_1372 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1374 = _T_1372 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1375 = _T_1372 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1376 = regs_6_15 + regs_6_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1696 = {{1'd0}, regs_6_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1377 = _T_1376 + _GEN_1696; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1697 = {{2'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1378 = _T_1377 + _GEN_1697; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1698 = {{3'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1379 = _T_1378 + _GEN_1698; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1699 = {{4'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1380 = _T_1379 + _GEN_1699; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1700 = {{5'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1381 = _T_1380 + _GEN_1700; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1701 = {{6'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1382 = _T_1381 + _GEN_1701; // @[Conwaylife.scala 31:34]
  wire  _T_1383 = _T_1382 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1384 = _T_1382 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1385 = _T_1382 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1386 = regs_6_0 + regs_6_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1702 = {{1'd0}, regs_6_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1387 = _T_1386 + _GEN_1702; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1703 = {{2'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1388 = _T_1387 + _GEN_1703; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1704 = {{3'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1389 = _T_1388 + _GEN_1704; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1705 = {{4'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1390 = _T_1389 + _GEN_1705; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1706 = {{5'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1391 = _T_1390 + _GEN_1706; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1707 = {{6'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1392 = _T_1391 + _GEN_1707; // @[Conwaylife.scala 31:34]
  wire  _T_1393 = _T_1392 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1394 = _T_1392 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1395 = _T_1392 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1396 = regs_6_1 + regs_6_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1708 = {{1'd0}, regs_6_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1397 = _T_1396 + _GEN_1708; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1709 = {{2'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1398 = _T_1397 + _GEN_1709; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1710 = {{3'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1399 = _T_1398 + _GEN_1710; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1711 = {{4'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1400 = _T_1399 + _GEN_1711; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1712 = {{5'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1401 = _T_1400 + _GEN_1712; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1713 = {{6'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1402 = _T_1401 + _GEN_1713; // @[Conwaylife.scala 31:34]
  wire  _T_1403 = _T_1402 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1404 = _T_1402 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1405 = _T_1402 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1406 = regs_6_2 + regs_6_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1714 = {{1'd0}, regs_6_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1407 = _T_1406 + _GEN_1714; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1715 = {{2'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1408 = _T_1407 + _GEN_1715; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1716 = {{3'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1409 = _T_1408 + _GEN_1716; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1717 = {{4'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1410 = _T_1409 + _GEN_1717; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1718 = {{5'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1411 = _T_1410 + _GEN_1718; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1719 = {{6'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1412 = _T_1411 + _GEN_1719; // @[Conwaylife.scala 31:34]
  wire  _T_1413 = _T_1412 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1414 = _T_1412 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1415 = _T_1412 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1416 = regs_6_3 + regs_6_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1720 = {{1'd0}, regs_6_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1417 = _T_1416 + _GEN_1720; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1721 = {{2'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1418 = _T_1417 + _GEN_1721; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1722 = {{3'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1419 = _T_1418 + _GEN_1722; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1723 = {{4'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1420 = _T_1419 + _GEN_1723; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1724 = {{5'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1421 = _T_1420 + _GEN_1724; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1725 = {{6'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1422 = _T_1421 + _GEN_1725; // @[Conwaylife.scala 31:34]
  wire  _T_1423 = _T_1422 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1424 = _T_1422 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1425 = _T_1422 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1426 = regs_6_4 + regs_6_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1726 = {{1'd0}, regs_6_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1427 = _T_1426 + _GEN_1726; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1727 = {{2'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1428 = _T_1427 + _GEN_1727; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1728 = {{3'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1429 = _T_1428 + _GEN_1728; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1729 = {{4'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1430 = _T_1429 + _GEN_1729; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1730 = {{5'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1431 = _T_1430 + _GEN_1730; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1731 = {{6'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1432 = _T_1431 + _GEN_1731; // @[Conwaylife.scala 31:34]
  wire  _T_1433 = _T_1432 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1434 = _T_1432 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1435 = _T_1432 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1436 = regs_6_5 + regs_6_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1732 = {{1'd0}, regs_6_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1437 = _T_1436 + _GEN_1732; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1733 = {{2'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1438 = _T_1437 + _GEN_1733; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1734 = {{3'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1439 = _T_1438 + _GEN_1734; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1735 = {{4'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1440 = _T_1439 + _GEN_1735; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1736 = {{5'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1441 = _T_1440 + _GEN_1736; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1737 = {{6'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1442 = _T_1441 + _GEN_1737; // @[Conwaylife.scala 31:34]
  wire  _T_1443 = _T_1442 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1444 = _T_1442 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1445 = _T_1442 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1446 = regs_6_6 + regs_6_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1738 = {{1'd0}, regs_6_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1447 = _T_1446 + _GEN_1738; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1739 = {{2'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1448 = _T_1447 + _GEN_1739; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1740 = {{3'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1449 = _T_1448 + _GEN_1740; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1741 = {{4'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1450 = _T_1449 + _GEN_1741; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1742 = {{5'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1451 = _T_1450 + _GEN_1742; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1743 = {{6'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1452 = _T_1451 + _GEN_1743; // @[Conwaylife.scala 31:34]
  wire  _T_1453 = _T_1452 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1454 = _T_1452 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1455 = _T_1452 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1456 = regs_6_7 + regs_6_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1744 = {{1'd0}, regs_6_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1457 = _T_1456 + _GEN_1744; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1745 = {{2'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1458 = _T_1457 + _GEN_1745; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1746 = {{3'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1459 = _T_1458 + _GEN_1746; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1747 = {{4'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1460 = _T_1459 + _GEN_1747; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1748 = {{5'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1461 = _T_1460 + _GEN_1748; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1749 = {{6'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1462 = _T_1461 + _GEN_1749; // @[Conwaylife.scala 31:34]
  wire  _T_1463 = _T_1462 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1464 = _T_1462 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1465 = _T_1462 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1466 = regs_6_8 + regs_6_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1750 = {{1'd0}, regs_6_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1467 = _T_1466 + _GEN_1750; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1751 = {{2'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1468 = _T_1467 + _GEN_1751; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1752 = {{3'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1469 = _T_1468 + _GEN_1752; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1753 = {{4'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1470 = _T_1469 + _GEN_1753; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1754 = {{5'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1471 = _T_1470 + _GEN_1754; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1755 = {{6'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1472 = _T_1471 + _GEN_1755; // @[Conwaylife.scala 31:34]
  wire  _T_1473 = _T_1472 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1474 = _T_1472 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1475 = _T_1472 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1476 = regs_6_9 + regs_6_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1756 = {{1'd0}, regs_6_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1477 = _T_1476 + _GEN_1756; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1757 = {{2'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1478 = _T_1477 + _GEN_1757; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1758 = {{3'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1479 = _T_1478 + _GEN_1758; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1759 = {{4'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1480 = _T_1479 + _GEN_1759; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1760 = {{5'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1481 = _T_1480 + _GEN_1760; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1761 = {{6'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1482 = _T_1481 + _GEN_1761; // @[Conwaylife.scala 31:34]
  wire  _T_1483 = _T_1482 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1484 = _T_1482 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1485 = _T_1482 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1486 = regs_6_10 + regs_6_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1762 = {{1'd0}, regs_6_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1487 = _T_1486 + _GEN_1762; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1763 = {{2'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1488 = _T_1487 + _GEN_1763; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1764 = {{3'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1489 = _T_1488 + _GEN_1764; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1765 = {{4'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1490 = _T_1489 + _GEN_1765; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1766 = {{5'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1491 = _T_1490 + _GEN_1766; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1767 = {{6'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1492 = _T_1491 + _GEN_1767; // @[Conwaylife.scala 31:34]
  wire  _T_1493 = _T_1492 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1494 = _T_1492 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1495 = _T_1492 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1496 = regs_6_11 + regs_6_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1768 = {{1'd0}, regs_6_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1497 = _T_1496 + _GEN_1768; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1769 = {{2'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1498 = _T_1497 + _GEN_1769; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1770 = {{3'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1499 = _T_1498 + _GEN_1770; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1771 = {{4'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1500 = _T_1499 + _GEN_1771; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1772 = {{5'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1501 = _T_1500 + _GEN_1772; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1773 = {{6'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1502 = _T_1501 + _GEN_1773; // @[Conwaylife.scala 31:34]
  wire  _T_1503 = _T_1502 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1504 = _T_1502 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1505 = _T_1502 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1506 = regs_6_12 + regs_6_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1774 = {{1'd0}, regs_6_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1507 = _T_1506 + _GEN_1774; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1775 = {{2'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1508 = _T_1507 + _GEN_1775; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1776 = {{3'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1509 = _T_1508 + _GEN_1776; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1777 = {{4'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1510 = _T_1509 + _GEN_1777; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1778 = {{5'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1511 = _T_1510 + _GEN_1778; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1779 = {{6'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1512 = _T_1511 + _GEN_1779; // @[Conwaylife.scala 31:34]
  wire  _T_1513 = _T_1512 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1514 = _T_1512 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1515 = _T_1512 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1516 = regs_6_13 + regs_6_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1780 = {{1'd0}, regs_6_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1517 = _T_1516 + _GEN_1780; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1781 = {{2'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1518 = _T_1517 + _GEN_1781; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1782 = {{3'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1519 = _T_1518 + _GEN_1782; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1783 = {{4'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1520 = _T_1519 + _GEN_1783; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1784 = {{5'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1521 = _T_1520 + _GEN_1784; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1785 = {{6'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1522 = _T_1521 + _GEN_1785; // @[Conwaylife.scala 31:34]
  wire  _T_1523 = _T_1522 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1524 = _T_1522 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1525 = _T_1522 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1526 = regs_6_14 + regs_6_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1786 = {{1'd0}, regs_6_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1527 = _T_1526 + _GEN_1786; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1787 = {{2'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1528 = _T_1527 + _GEN_1787; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1788 = {{3'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1529 = _T_1528 + _GEN_1788; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1789 = {{4'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1530 = _T_1529 + _GEN_1789; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1790 = {{5'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1531 = _T_1530 + _GEN_1790; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1791 = {{6'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1532 = _T_1531 + _GEN_1791; // @[Conwaylife.scala 31:34]
  wire  _T_1533 = _T_1532 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1534 = _T_1532 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1535 = _T_1532 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1536 = regs_7_15 + regs_7_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1792 = {{1'd0}, regs_7_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1537 = _T_1536 + _GEN_1792; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1793 = {{2'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1538 = _T_1537 + _GEN_1793; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1794 = {{3'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1539 = _T_1538 + _GEN_1794; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1795 = {{4'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1540 = _T_1539 + _GEN_1795; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1796 = {{5'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1541 = _T_1540 + _GEN_1796; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1797 = {{6'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1542 = _T_1541 + _GEN_1797; // @[Conwaylife.scala 31:34]
  wire  _T_1543 = _T_1542 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1544 = _T_1542 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1545 = _T_1542 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1546 = regs_7_0 + regs_7_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1798 = {{1'd0}, regs_7_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1547 = _T_1546 + _GEN_1798; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1799 = {{2'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1548 = _T_1547 + _GEN_1799; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1800 = {{3'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1549 = _T_1548 + _GEN_1800; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1801 = {{4'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1550 = _T_1549 + _GEN_1801; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1802 = {{5'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1551 = _T_1550 + _GEN_1802; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1803 = {{6'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1552 = _T_1551 + _GEN_1803; // @[Conwaylife.scala 31:34]
  wire  _T_1553 = _T_1552 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1554 = _T_1552 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1555 = _T_1552 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1556 = regs_7_1 + regs_7_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1804 = {{1'd0}, regs_7_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1557 = _T_1556 + _GEN_1804; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1805 = {{2'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1558 = _T_1557 + _GEN_1805; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1806 = {{3'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1559 = _T_1558 + _GEN_1806; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1807 = {{4'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1560 = _T_1559 + _GEN_1807; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1808 = {{5'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1561 = _T_1560 + _GEN_1808; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1809 = {{6'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1562 = _T_1561 + _GEN_1809; // @[Conwaylife.scala 31:34]
  wire  _T_1563 = _T_1562 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1564 = _T_1562 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1565 = _T_1562 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1566 = regs_7_2 + regs_7_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1810 = {{1'd0}, regs_7_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1567 = _T_1566 + _GEN_1810; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1811 = {{2'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1568 = _T_1567 + _GEN_1811; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1812 = {{3'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1569 = _T_1568 + _GEN_1812; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1813 = {{4'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1570 = _T_1569 + _GEN_1813; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1814 = {{5'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1571 = _T_1570 + _GEN_1814; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1815 = {{6'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1572 = _T_1571 + _GEN_1815; // @[Conwaylife.scala 31:34]
  wire  _T_1573 = _T_1572 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1574 = _T_1572 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1575 = _T_1572 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1576 = regs_7_3 + regs_7_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1816 = {{1'd0}, regs_7_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1577 = _T_1576 + _GEN_1816; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1817 = {{2'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1578 = _T_1577 + _GEN_1817; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1818 = {{3'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1579 = _T_1578 + _GEN_1818; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1819 = {{4'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1580 = _T_1579 + _GEN_1819; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1820 = {{5'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1581 = _T_1580 + _GEN_1820; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1821 = {{6'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1582 = _T_1581 + _GEN_1821; // @[Conwaylife.scala 31:34]
  wire  _T_1583 = _T_1582 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1584 = _T_1582 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1585 = _T_1582 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1586 = regs_7_4 + regs_7_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1822 = {{1'd0}, regs_7_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1587 = _T_1586 + _GEN_1822; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1823 = {{2'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1588 = _T_1587 + _GEN_1823; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1824 = {{3'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1589 = _T_1588 + _GEN_1824; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1825 = {{4'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1590 = _T_1589 + _GEN_1825; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1826 = {{5'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1591 = _T_1590 + _GEN_1826; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1827 = {{6'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1592 = _T_1591 + _GEN_1827; // @[Conwaylife.scala 31:34]
  wire  _T_1593 = _T_1592 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1594 = _T_1592 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1595 = _T_1592 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1596 = regs_7_5 + regs_7_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1828 = {{1'd0}, regs_7_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1597 = _T_1596 + _GEN_1828; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1829 = {{2'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1598 = _T_1597 + _GEN_1829; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1830 = {{3'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1599 = _T_1598 + _GEN_1830; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1831 = {{4'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1600 = _T_1599 + _GEN_1831; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1832 = {{5'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1601 = _T_1600 + _GEN_1832; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1833 = {{6'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1602 = _T_1601 + _GEN_1833; // @[Conwaylife.scala 31:34]
  wire  _T_1603 = _T_1602 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1604 = _T_1602 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1605 = _T_1602 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1606 = regs_7_6 + regs_7_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1834 = {{1'd0}, regs_7_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1607 = _T_1606 + _GEN_1834; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1835 = {{2'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1608 = _T_1607 + _GEN_1835; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1836 = {{3'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1609 = _T_1608 + _GEN_1836; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1837 = {{4'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1610 = _T_1609 + _GEN_1837; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1838 = {{5'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1611 = _T_1610 + _GEN_1838; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1839 = {{6'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1612 = _T_1611 + _GEN_1839; // @[Conwaylife.scala 31:34]
  wire  _T_1613 = _T_1612 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1614 = _T_1612 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1615 = _T_1612 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1616 = regs_7_7 + regs_7_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1840 = {{1'd0}, regs_7_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1617 = _T_1616 + _GEN_1840; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1841 = {{2'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1618 = _T_1617 + _GEN_1841; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1842 = {{3'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1619 = _T_1618 + _GEN_1842; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1843 = {{4'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1620 = _T_1619 + _GEN_1843; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1844 = {{5'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1621 = _T_1620 + _GEN_1844; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1845 = {{6'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1622 = _T_1621 + _GEN_1845; // @[Conwaylife.scala 31:34]
  wire  _T_1623 = _T_1622 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1624 = _T_1622 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1625 = _T_1622 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1626 = regs_7_8 + regs_7_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1846 = {{1'd0}, regs_7_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1627 = _T_1626 + _GEN_1846; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1847 = {{2'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1628 = _T_1627 + _GEN_1847; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1848 = {{3'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1629 = _T_1628 + _GEN_1848; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1849 = {{4'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1630 = _T_1629 + _GEN_1849; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1850 = {{5'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1631 = _T_1630 + _GEN_1850; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1851 = {{6'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1632 = _T_1631 + _GEN_1851; // @[Conwaylife.scala 31:34]
  wire  _T_1633 = _T_1632 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1634 = _T_1632 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1635 = _T_1632 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1636 = regs_7_9 + regs_7_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1852 = {{1'd0}, regs_7_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1637 = _T_1636 + _GEN_1852; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1853 = {{2'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1638 = _T_1637 + _GEN_1853; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1854 = {{3'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1639 = _T_1638 + _GEN_1854; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1855 = {{4'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1640 = _T_1639 + _GEN_1855; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1856 = {{5'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1641 = _T_1640 + _GEN_1856; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1857 = {{6'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1642 = _T_1641 + _GEN_1857; // @[Conwaylife.scala 31:34]
  wire  _T_1643 = _T_1642 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1644 = _T_1642 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1645 = _T_1642 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1646 = regs_7_10 + regs_7_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1858 = {{1'd0}, regs_7_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1647 = _T_1646 + _GEN_1858; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1859 = {{2'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1648 = _T_1647 + _GEN_1859; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1860 = {{3'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1649 = _T_1648 + _GEN_1860; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1861 = {{4'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1650 = _T_1649 + _GEN_1861; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1862 = {{5'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1651 = _T_1650 + _GEN_1862; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1863 = {{6'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1652 = _T_1651 + _GEN_1863; // @[Conwaylife.scala 31:34]
  wire  _T_1653 = _T_1652 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1654 = _T_1652 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1655 = _T_1652 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1656 = regs_7_11 + regs_7_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1864 = {{1'd0}, regs_7_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1657 = _T_1656 + _GEN_1864; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1865 = {{2'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1658 = _T_1657 + _GEN_1865; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1866 = {{3'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1659 = _T_1658 + _GEN_1866; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1867 = {{4'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1660 = _T_1659 + _GEN_1867; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1868 = {{5'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1661 = _T_1660 + _GEN_1868; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1869 = {{6'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1662 = _T_1661 + _GEN_1869; // @[Conwaylife.scala 31:34]
  wire  _T_1663 = _T_1662 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1664 = _T_1662 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1665 = _T_1662 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1666 = regs_7_12 + regs_7_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1870 = {{1'd0}, regs_7_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1667 = _T_1666 + _GEN_1870; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1871 = {{2'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1668 = _T_1667 + _GEN_1871; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1872 = {{3'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1669 = _T_1668 + _GEN_1872; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1873 = {{4'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1670 = _T_1669 + _GEN_1873; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1874 = {{5'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1671 = _T_1670 + _GEN_1874; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1875 = {{6'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1672 = _T_1671 + _GEN_1875; // @[Conwaylife.scala 31:34]
  wire  _T_1673 = _T_1672 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1674 = _T_1672 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1675 = _T_1672 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1676 = regs_7_13 + regs_7_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1876 = {{1'd0}, regs_7_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1677 = _T_1676 + _GEN_1876; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1877 = {{2'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1678 = _T_1677 + _GEN_1877; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1878 = {{3'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1679 = _T_1678 + _GEN_1878; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1879 = {{4'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1680 = _T_1679 + _GEN_1879; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1880 = {{5'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1681 = _T_1680 + _GEN_1880; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1881 = {{6'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1682 = _T_1681 + _GEN_1881; // @[Conwaylife.scala 31:34]
  wire  _T_1683 = _T_1682 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1684 = _T_1682 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1685 = _T_1682 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1686 = regs_7_14 + regs_7_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1882 = {{1'd0}, regs_7_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1687 = _T_1686 + _GEN_1882; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1883 = {{2'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1688 = _T_1687 + _GEN_1883; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1884 = {{3'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1689 = _T_1688 + _GEN_1884; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1885 = {{4'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1690 = _T_1689 + _GEN_1885; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1886 = {{5'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1691 = _T_1690 + _GEN_1886; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1887 = {{6'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1692 = _T_1691 + _GEN_1887; // @[Conwaylife.scala 31:34]
  wire  _T_1693 = _T_1692 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1694 = _T_1692 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1695 = _T_1692 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1696 = regs_8_15 + regs_8_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1888 = {{1'd0}, regs_8_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1697 = _T_1696 + _GEN_1888; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1889 = {{2'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1698 = _T_1697 + _GEN_1889; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1890 = {{3'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1699 = _T_1698 + _GEN_1890; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1891 = {{4'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1700 = _T_1699 + _GEN_1891; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1892 = {{5'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1701 = _T_1700 + _GEN_1892; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1893 = {{6'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1702 = _T_1701 + _GEN_1893; // @[Conwaylife.scala 31:34]
  wire  _T_1703 = _T_1702 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1704 = _T_1702 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1705 = _T_1702 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1706 = regs_8_0 + regs_8_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1894 = {{1'd0}, regs_8_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1707 = _T_1706 + _GEN_1894; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1895 = {{2'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1708 = _T_1707 + _GEN_1895; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1896 = {{3'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1709 = _T_1708 + _GEN_1896; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1897 = {{4'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1710 = _T_1709 + _GEN_1897; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1898 = {{5'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1711 = _T_1710 + _GEN_1898; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1899 = {{6'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1712 = _T_1711 + _GEN_1899; // @[Conwaylife.scala 31:34]
  wire  _T_1713 = _T_1712 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1714 = _T_1712 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1715 = _T_1712 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1716 = regs_8_1 + regs_8_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1900 = {{1'd0}, regs_8_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1717 = _T_1716 + _GEN_1900; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1901 = {{2'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1718 = _T_1717 + _GEN_1901; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1902 = {{3'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1719 = _T_1718 + _GEN_1902; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1903 = {{4'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1720 = _T_1719 + _GEN_1903; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1904 = {{5'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1721 = _T_1720 + _GEN_1904; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1905 = {{6'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1722 = _T_1721 + _GEN_1905; // @[Conwaylife.scala 31:34]
  wire  _T_1723 = _T_1722 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1724 = _T_1722 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1725 = _T_1722 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1726 = regs_8_2 + regs_8_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1906 = {{1'd0}, regs_8_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1727 = _T_1726 + _GEN_1906; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1907 = {{2'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1728 = _T_1727 + _GEN_1907; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1908 = {{3'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1729 = _T_1728 + _GEN_1908; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1909 = {{4'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1730 = _T_1729 + _GEN_1909; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1910 = {{5'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1731 = _T_1730 + _GEN_1910; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1911 = {{6'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1732 = _T_1731 + _GEN_1911; // @[Conwaylife.scala 31:34]
  wire  _T_1733 = _T_1732 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1734 = _T_1732 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1735 = _T_1732 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1736 = regs_8_3 + regs_8_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1912 = {{1'd0}, regs_8_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1737 = _T_1736 + _GEN_1912; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1913 = {{2'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1738 = _T_1737 + _GEN_1913; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1914 = {{3'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1739 = _T_1738 + _GEN_1914; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1915 = {{4'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1740 = _T_1739 + _GEN_1915; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1916 = {{5'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1741 = _T_1740 + _GEN_1916; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1917 = {{6'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1742 = _T_1741 + _GEN_1917; // @[Conwaylife.scala 31:34]
  wire  _T_1743 = _T_1742 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1744 = _T_1742 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1745 = _T_1742 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1746 = regs_8_4 + regs_8_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1918 = {{1'd0}, regs_8_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1747 = _T_1746 + _GEN_1918; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1919 = {{2'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1748 = _T_1747 + _GEN_1919; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1920 = {{3'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1749 = _T_1748 + _GEN_1920; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1921 = {{4'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1750 = _T_1749 + _GEN_1921; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1922 = {{5'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1751 = _T_1750 + _GEN_1922; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1923 = {{6'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1752 = _T_1751 + _GEN_1923; // @[Conwaylife.scala 31:34]
  wire  _T_1753 = _T_1752 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1754 = _T_1752 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1755 = _T_1752 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1756 = regs_8_5 + regs_8_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1924 = {{1'd0}, regs_8_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1757 = _T_1756 + _GEN_1924; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1925 = {{2'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1758 = _T_1757 + _GEN_1925; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1926 = {{3'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1759 = _T_1758 + _GEN_1926; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1927 = {{4'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1760 = _T_1759 + _GEN_1927; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1928 = {{5'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1761 = _T_1760 + _GEN_1928; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1929 = {{6'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1762 = _T_1761 + _GEN_1929; // @[Conwaylife.scala 31:34]
  wire  _T_1763 = _T_1762 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1764 = _T_1762 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1765 = _T_1762 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1766 = regs_8_6 + regs_8_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1930 = {{1'd0}, regs_8_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1767 = _T_1766 + _GEN_1930; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1931 = {{2'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1768 = _T_1767 + _GEN_1931; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1932 = {{3'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1769 = _T_1768 + _GEN_1932; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1933 = {{4'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1770 = _T_1769 + _GEN_1933; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1934 = {{5'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1771 = _T_1770 + _GEN_1934; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1935 = {{6'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1772 = _T_1771 + _GEN_1935; // @[Conwaylife.scala 31:34]
  wire  _T_1773 = _T_1772 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1774 = _T_1772 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1775 = _T_1772 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1776 = regs_8_7 + regs_8_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1936 = {{1'd0}, regs_8_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1777 = _T_1776 + _GEN_1936; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1937 = {{2'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1778 = _T_1777 + _GEN_1937; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1938 = {{3'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1779 = _T_1778 + _GEN_1938; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1939 = {{4'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1780 = _T_1779 + _GEN_1939; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1940 = {{5'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1781 = _T_1780 + _GEN_1940; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1941 = {{6'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1782 = _T_1781 + _GEN_1941; // @[Conwaylife.scala 31:34]
  wire  _T_1783 = _T_1782 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1784 = _T_1782 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1785 = _T_1782 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1786 = regs_8_8 + regs_8_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1942 = {{1'd0}, regs_8_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1787 = _T_1786 + _GEN_1942; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1943 = {{2'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1788 = _T_1787 + _GEN_1943; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1944 = {{3'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1789 = _T_1788 + _GEN_1944; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1945 = {{4'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1790 = _T_1789 + _GEN_1945; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1946 = {{5'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1791 = _T_1790 + _GEN_1946; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1947 = {{6'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1792 = _T_1791 + _GEN_1947; // @[Conwaylife.scala 31:34]
  wire  _T_1793 = _T_1792 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1794 = _T_1792 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1795 = _T_1792 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1796 = regs_8_9 + regs_8_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1948 = {{1'd0}, regs_8_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1797 = _T_1796 + _GEN_1948; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1949 = {{2'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1798 = _T_1797 + _GEN_1949; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1950 = {{3'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1799 = _T_1798 + _GEN_1950; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1951 = {{4'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1800 = _T_1799 + _GEN_1951; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1952 = {{5'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1801 = _T_1800 + _GEN_1952; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1953 = {{6'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1802 = _T_1801 + _GEN_1953; // @[Conwaylife.scala 31:34]
  wire  _T_1803 = _T_1802 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1804 = _T_1802 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1805 = _T_1802 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1806 = regs_8_10 + regs_8_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1954 = {{1'd0}, regs_8_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1807 = _T_1806 + _GEN_1954; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1955 = {{2'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1808 = _T_1807 + _GEN_1955; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1956 = {{3'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1809 = _T_1808 + _GEN_1956; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1957 = {{4'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1810 = _T_1809 + _GEN_1957; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1958 = {{5'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1811 = _T_1810 + _GEN_1958; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1959 = {{6'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1812 = _T_1811 + _GEN_1959; // @[Conwaylife.scala 31:34]
  wire  _T_1813 = _T_1812 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1814 = _T_1812 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1815 = _T_1812 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1816 = regs_8_11 + regs_8_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1960 = {{1'd0}, regs_8_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1817 = _T_1816 + _GEN_1960; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1961 = {{2'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1818 = _T_1817 + _GEN_1961; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1962 = {{3'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1819 = _T_1818 + _GEN_1962; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1963 = {{4'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1820 = _T_1819 + _GEN_1963; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1964 = {{5'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1821 = _T_1820 + _GEN_1964; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1965 = {{6'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1822 = _T_1821 + _GEN_1965; // @[Conwaylife.scala 31:34]
  wire  _T_1823 = _T_1822 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1824 = _T_1822 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1825 = _T_1822 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1826 = regs_8_12 + regs_8_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1966 = {{1'd0}, regs_8_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1827 = _T_1826 + _GEN_1966; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1967 = {{2'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1828 = _T_1827 + _GEN_1967; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1968 = {{3'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1829 = _T_1828 + _GEN_1968; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1969 = {{4'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1830 = _T_1829 + _GEN_1969; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1970 = {{5'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1831 = _T_1830 + _GEN_1970; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1971 = {{6'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1832 = _T_1831 + _GEN_1971; // @[Conwaylife.scala 31:34]
  wire  _T_1833 = _T_1832 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1834 = _T_1832 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1835 = _T_1832 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1836 = regs_8_13 + regs_8_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1972 = {{1'd0}, regs_8_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1837 = _T_1836 + _GEN_1972; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1973 = {{2'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1838 = _T_1837 + _GEN_1973; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1974 = {{3'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1839 = _T_1838 + _GEN_1974; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1975 = {{4'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1840 = _T_1839 + _GEN_1975; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1976 = {{5'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1841 = _T_1840 + _GEN_1976; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1977 = {{6'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1842 = _T_1841 + _GEN_1977; // @[Conwaylife.scala 31:34]
  wire  _T_1843 = _T_1842 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1844 = _T_1842 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1845 = _T_1842 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1846 = regs_8_14 + regs_8_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1978 = {{1'd0}, regs_8_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1847 = _T_1846 + _GEN_1978; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1979 = {{2'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1848 = _T_1847 + _GEN_1979; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1980 = {{3'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1849 = _T_1848 + _GEN_1980; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1981 = {{4'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1850 = _T_1849 + _GEN_1981; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1982 = {{5'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1851 = _T_1850 + _GEN_1982; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1983 = {{6'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1852 = _T_1851 + _GEN_1983; // @[Conwaylife.scala 31:34]
  wire  _T_1853 = _T_1852 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1854 = _T_1852 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1855 = _T_1852 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1856 = regs_9_15 + regs_9_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1984 = {{1'd0}, regs_9_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1857 = _T_1856 + _GEN_1984; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1985 = {{2'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1858 = _T_1857 + _GEN_1985; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1986 = {{3'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1859 = _T_1858 + _GEN_1986; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1987 = {{4'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1860 = _T_1859 + _GEN_1987; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1988 = {{5'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1861 = _T_1860 + _GEN_1988; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1989 = {{6'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1862 = _T_1861 + _GEN_1989; // @[Conwaylife.scala 31:34]
  wire  _T_1863 = _T_1862 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1864 = _T_1862 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1865 = _T_1862 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1866 = regs_9_0 + regs_9_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1990 = {{1'd0}, regs_9_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1867 = _T_1866 + _GEN_1990; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1991 = {{2'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1868 = _T_1867 + _GEN_1991; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1992 = {{3'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1869 = _T_1868 + _GEN_1992; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1993 = {{4'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1870 = _T_1869 + _GEN_1993; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_1994 = {{5'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1871 = _T_1870 + _GEN_1994; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_1995 = {{6'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1872 = _T_1871 + _GEN_1995; // @[Conwaylife.scala 31:34]
  wire  _T_1873 = _T_1872 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1874 = _T_1872 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1875 = _T_1872 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1876 = regs_9_1 + regs_9_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_1996 = {{1'd0}, regs_9_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1877 = _T_1876 + _GEN_1996; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_1997 = {{2'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1878 = _T_1877 + _GEN_1997; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_1998 = {{3'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1879 = _T_1878 + _GEN_1998; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_1999 = {{4'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1880 = _T_1879 + _GEN_1999; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2000 = {{5'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1881 = _T_1880 + _GEN_2000; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2001 = {{6'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1882 = _T_1881 + _GEN_2001; // @[Conwaylife.scala 31:34]
  wire  _T_1883 = _T_1882 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1884 = _T_1882 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1885 = _T_1882 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1886 = regs_9_2 + regs_9_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2002 = {{1'd0}, regs_9_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1887 = _T_1886 + _GEN_2002; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2003 = {{2'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1888 = _T_1887 + _GEN_2003; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2004 = {{3'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1889 = _T_1888 + _GEN_2004; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2005 = {{4'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1890 = _T_1889 + _GEN_2005; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2006 = {{5'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1891 = _T_1890 + _GEN_2006; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2007 = {{6'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1892 = _T_1891 + _GEN_2007; // @[Conwaylife.scala 31:34]
  wire  _T_1893 = _T_1892 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1894 = _T_1892 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1895 = _T_1892 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1896 = regs_9_3 + regs_9_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2008 = {{1'd0}, regs_9_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1897 = _T_1896 + _GEN_2008; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2009 = {{2'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1898 = _T_1897 + _GEN_2009; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2010 = {{3'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1899 = _T_1898 + _GEN_2010; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2011 = {{4'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1900 = _T_1899 + _GEN_2011; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2012 = {{5'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1901 = _T_1900 + _GEN_2012; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2013 = {{6'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1902 = _T_1901 + _GEN_2013; // @[Conwaylife.scala 31:34]
  wire  _T_1903 = _T_1902 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1904 = _T_1902 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1905 = _T_1902 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1906 = regs_9_4 + regs_9_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2014 = {{1'd0}, regs_9_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1907 = _T_1906 + _GEN_2014; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2015 = {{2'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1908 = _T_1907 + _GEN_2015; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2016 = {{3'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1909 = _T_1908 + _GEN_2016; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2017 = {{4'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1910 = _T_1909 + _GEN_2017; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2018 = {{5'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1911 = _T_1910 + _GEN_2018; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2019 = {{6'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1912 = _T_1911 + _GEN_2019; // @[Conwaylife.scala 31:34]
  wire  _T_1913 = _T_1912 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1914 = _T_1912 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1915 = _T_1912 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1916 = regs_9_5 + regs_9_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2020 = {{1'd0}, regs_9_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1917 = _T_1916 + _GEN_2020; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2021 = {{2'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1918 = _T_1917 + _GEN_2021; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2022 = {{3'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1919 = _T_1918 + _GEN_2022; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2023 = {{4'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1920 = _T_1919 + _GEN_2023; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2024 = {{5'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1921 = _T_1920 + _GEN_2024; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2025 = {{6'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1922 = _T_1921 + _GEN_2025; // @[Conwaylife.scala 31:34]
  wire  _T_1923 = _T_1922 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1924 = _T_1922 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1925 = _T_1922 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1926 = regs_9_6 + regs_9_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2026 = {{1'd0}, regs_9_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1927 = _T_1926 + _GEN_2026; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2027 = {{2'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1928 = _T_1927 + _GEN_2027; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2028 = {{3'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1929 = _T_1928 + _GEN_2028; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2029 = {{4'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1930 = _T_1929 + _GEN_2029; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2030 = {{5'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1931 = _T_1930 + _GEN_2030; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2031 = {{6'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1932 = _T_1931 + _GEN_2031; // @[Conwaylife.scala 31:34]
  wire  _T_1933 = _T_1932 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1934 = _T_1932 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1935 = _T_1932 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1936 = regs_9_7 + regs_9_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2032 = {{1'd0}, regs_9_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1937 = _T_1936 + _GEN_2032; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2033 = {{2'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1938 = _T_1937 + _GEN_2033; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2034 = {{3'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1939 = _T_1938 + _GEN_2034; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2035 = {{4'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1940 = _T_1939 + _GEN_2035; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2036 = {{5'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1941 = _T_1940 + _GEN_2036; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2037 = {{6'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1942 = _T_1941 + _GEN_2037; // @[Conwaylife.scala 31:34]
  wire  _T_1943 = _T_1942 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1944 = _T_1942 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1945 = _T_1942 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1946 = regs_9_8 + regs_9_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2038 = {{1'd0}, regs_9_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1947 = _T_1946 + _GEN_2038; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2039 = {{2'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1948 = _T_1947 + _GEN_2039; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2040 = {{3'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1949 = _T_1948 + _GEN_2040; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2041 = {{4'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1950 = _T_1949 + _GEN_2041; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2042 = {{5'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1951 = _T_1950 + _GEN_2042; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2043 = {{6'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1952 = _T_1951 + _GEN_2043; // @[Conwaylife.scala 31:34]
  wire  _T_1953 = _T_1952 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1954 = _T_1952 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1955 = _T_1952 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1956 = regs_9_9 + regs_9_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2044 = {{1'd0}, regs_9_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1957 = _T_1956 + _GEN_2044; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2045 = {{2'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1958 = _T_1957 + _GEN_2045; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2046 = {{3'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1959 = _T_1958 + _GEN_2046; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2047 = {{4'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1960 = _T_1959 + _GEN_2047; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2048 = {{5'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1961 = _T_1960 + _GEN_2048; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2049 = {{6'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1962 = _T_1961 + _GEN_2049; // @[Conwaylife.scala 31:34]
  wire  _T_1963 = _T_1962 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1964 = _T_1962 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1965 = _T_1962 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1966 = regs_9_10 + regs_9_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2050 = {{1'd0}, regs_9_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1967 = _T_1966 + _GEN_2050; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2051 = {{2'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1968 = _T_1967 + _GEN_2051; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2052 = {{3'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1969 = _T_1968 + _GEN_2052; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2053 = {{4'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1970 = _T_1969 + _GEN_2053; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2054 = {{5'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1971 = _T_1970 + _GEN_2054; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2055 = {{6'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1972 = _T_1971 + _GEN_2055; // @[Conwaylife.scala 31:34]
  wire  _T_1973 = _T_1972 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1974 = _T_1972 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1975 = _T_1972 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1976 = regs_9_11 + regs_9_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2056 = {{1'd0}, regs_9_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1977 = _T_1976 + _GEN_2056; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2057 = {{2'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1978 = _T_1977 + _GEN_2057; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2058 = {{3'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1979 = _T_1978 + _GEN_2058; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2059 = {{4'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1980 = _T_1979 + _GEN_2059; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2060 = {{5'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1981 = _T_1980 + _GEN_2060; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2061 = {{6'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1982 = _T_1981 + _GEN_2061; // @[Conwaylife.scala 31:34]
  wire  _T_1983 = _T_1982 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1984 = _T_1982 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1985 = _T_1982 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1986 = regs_9_12 + regs_9_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2062 = {{1'd0}, regs_9_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1987 = _T_1986 + _GEN_2062; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2063 = {{2'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1988 = _T_1987 + _GEN_2063; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2064 = {{3'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1989 = _T_1988 + _GEN_2064; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2065 = {{4'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_1990 = _T_1989 + _GEN_2065; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2066 = {{5'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_1991 = _T_1990 + _GEN_2066; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2067 = {{6'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_1992 = _T_1991 + _GEN_2067; // @[Conwaylife.scala 31:34]
  wire  _T_1993 = _T_1992 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_1994 = _T_1992 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_1995 = _T_1992 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_1996 = regs_9_13 + regs_9_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2068 = {{1'd0}, regs_9_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_1997 = _T_1996 + _GEN_2068; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2069 = {{2'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_1998 = _T_1997 + _GEN_2069; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2070 = {{3'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_1999 = _T_1998 + _GEN_2070; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2071 = {{4'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2000 = _T_1999 + _GEN_2071; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2072 = {{5'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2001 = _T_2000 + _GEN_2072; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2073 = {{6'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2002 = _T_2001 + _GEN_2073; // @[Conwaylife.scala 31:34]
  wire  _T_2003 = _T_2002 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2004 = _T_2002 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2005 = _T_2002 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2006 = regs_9_14 + regs_9_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2074 = {{1'd0}, regs_9_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2007 = _T_2006 + _GEN_2074; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2075 = {{2'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2008 = _T_2007 + _GEN_2075; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2076 = {{3'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2009 = _T_2008 + _GEN_2076; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2077 = {{4'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2010 = _T_2009 + _GEN_2077; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2078 = {{5'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2011 = _T_2010 + _GEN_2078; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2079 = {{6'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2012 = _T_2011 + _GEN_2079; // @[Conwaylife.scala 31:34]
  wire  _T_2013 = _T_2012 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2014 = _T_2012 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2015 = _T_2012 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2016 = regs_10_15 + regs_10_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2080 = {{1'd0}, regs_10_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2017 = _T_2016 + _GEN_2080; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2081 = {{2'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2018 = _T_2017 + _GEN_2081; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2082 = {{3'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2019 = _T_2018 + _GEN_2082; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2083 = {{4'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2020 = _T_2019 + _GEN_2083; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2084 = {{5'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2021 = _T_2020 + _GEN_2084; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2085 = {{6'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2022 = _T_2021 + _GEN_2085; // @[Conwaylife.scala 31:34]
  wire  _T_2023 = _T_2022 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2024 = _T_2022 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2025 = _T_2022 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2026 = regs_10_0 + regs_10_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2086 = {{1'd0}, regs_10_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2027 = _T_2026 + _GEN_2086; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2087 = {{2'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2028 = _T_2027 + _GEN_2087; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2088 = {{3'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2029 = _T_2028 + _GEN_2088; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2089 = {{4'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2030 = _T_2029 + _GEN_2089; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2090 = {{5'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2031 = _T_2030 + _GEN_2090; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2091 = {{6'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2032 = _T_2031 + _GEN_2091; // @[Conwaylife.scala 31:34]
  wire  _T_2033 = _T_2032 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2034 = _T_2032 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2035 = _T_2032 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2036 = regs_10_1 + regs_10_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2092 = {{1'd0}, regs_10_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2037 = _T_2036 + _GEN_2092; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2093 = {{2'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2038 = _T_2037 + _GEN_2093; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2094 = {{3'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2039 = _T_2038 + _GEN_2094; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2095 = {{4'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2040 = _T_2039 + _GEN_2095; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2096 = {{5'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2041 = _T_2040 + _GEN_2096; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2097 = {{6'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2042 = _T_2041 + _GEN_2097; // @[Conwaylife.scala 31:34]
  wire  _T_2043 = _T_2042 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2044 = _T_2042 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2045 = _T_2042 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2046 = regs_10_2 + regs_10_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2098 = {{1'd0}, regs_10_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2047 = _T_2046 + _GEN_2098; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2099 = {{2'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2048 = _T_2047 + _GEN_2099; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2100 = {{3'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2049 = _T_2048 + _GEN_2100; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2101 = {{4'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2050 = _T_2049 + _GEN_2101; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2102 = {{5'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2051 = _T_2050 + _GEN_2102; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2103 = {{6'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2052 = _T_2051 + _GEN_2103; // @[Conwaylife.scala 31:34]
  wire  _T_2053 = _T_2052 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2054 = _T_2052 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2055 = _T_2052 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2056 = regs_10_3 + regs_10_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2104 = {{1'd0}, regs_10_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2057 = _T_2056 + _GEN_2104; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2105 = {{2'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2058 = _T_2057 + _GEN_2105; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2106 = {{3'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2059 = _T_2058 + _GEN_2106; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2107 = {{4'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2060 = _T_2059 + _GEN_2107; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2108 = {{5'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2061 = _T_2060 + _GEN_2108; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2109 = {{6'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2062 = _T_2061 + _GEN_2109; // @[Conwaylife.scala 31:34]
  wire  _T_2063 = _T_2062 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2064 = _T_2062 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2065 = _T_2062 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2066 = regs_10_4 + regs_10_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2110 = {{1'd0}, regs_10_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2067 = _T_2066 + _GEN_2110; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2111 = {{2'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2068 = _T_2067 + _GEN_2111; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2112 = {{3'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2069 = _T_2068 + _GEN_2112; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2113 = {{4'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2070 = _T_2069 + _GEN_2113; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2114 = {{5'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2071 = _T_2070 + _GEN_2114; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2115 = {{6'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2072 = _T_2071 + _GEN_2115; // @[Conwaylife.scala 31:34]
  wire  _T_2073 = _T_2072 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2074 = _T_2072 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2075 = _T_2072 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2076 = regs_10_5 + regs_10_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2116 = {{1'd0}, regs_10_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2077 = _T_2076 + _GEN_2116; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2117 = {{2'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2078 = _T_2077 + _GEN_2117; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2118 = {{3'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2079 = _T_2078 + _GEN_2118; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2119 = {{4'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2080 = _T_2079 + _GEN_2119; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2120 = {{5'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2081 = _T_2080 + _GEN_2120; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2121 = {{6'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2082 = _T_2081 + _GEN_2121; // @[Conwaylife.scala 31:34]
  wire  _T_2083 = _T_2082 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2084 = _T_2082 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2085 = _T_2082 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2086 = regs_10_6 + regs_10_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2122 = {{1'd0}, regs_10_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2087 = _T_2086 + _GEN_2122; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2123 = {{2'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2088 = _T_2087 + _GEN_2123; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2124 = {{3'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2089 = _T_2088 + _GEN_2124; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2125 = {{4'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2090 = _T_2089 + _GEN_2125; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2126 = {{5'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2091 = _T_2090 + _GEN_2126; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2127 = {{6'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2092 = _T_2091 + _GEN_2127; // @[Conwaylife.scala 31:34]
  wire  _T_2093 = _T_2092 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2094 = _T_2092 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2095 = _T_2092 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2096 = regs_10_7 + regs_10_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2128 = {{1'd0}, regs_10_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2097 = _T_2096 + _GEN_2128; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2129 = {{2'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2098 = _T_2097 + _GEN_2129; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2130 = {{3'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2099 = _T_2098 + _GEN_2130; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2131 = {{4'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2100 = _T_2099 + _GEN_2131; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2132 = {{5'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2101 = _T_2100 + _GEN_2132; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2133 = {{6'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2102 = _T_2101 + _GEN_2133; // @[Conwaylife.scala 31:34]
  wire  _T_2103 = _T_2102 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2104 = _T_2102 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2105 = _T_2102 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2106 = regs_10_8 + regs_10_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2134 = {{1'd0}, regs_10_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2107 = _T_2106 + _GEN_2134; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2135 = {{2'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2108 = _T_2107 + _GEN_2135; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2136 = {{3'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2109 = _T_2108 + _GEN_2136; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2137 = {{4'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2110 = _T_2109 + _GEN_2137; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2138 = {{5'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2111 = _T_2110 + _GEN_2138; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2139 = {{6'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2112 = _T_2111 + _GEN_2139; // @[Conwaylife.scala 31:34]
  wire  _T_2113 = _T_2112 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2114 = _T_2112 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2115 = _T_2112 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2116 = regs_10_9 + regs_10_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2140 = {{1'd0}, regs_10_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2117 = _T_2116 + _GEN_2140; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2141 = {{2'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2118 = _T_2117 + _GEN_2141; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2142 = {{3'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2119 = _T_2118 + _GEN_2142; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2143 = {{4'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2120 = _T_2119 + _GEN_2143; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2144 = {{5'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2121 = _T_2120 + _GEN_2144; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2145 = {{6'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2122 = _T_2121 + _GEN_2145; // @[Conwaylife.scala 31:34]
  wire  _T_2123 = _T_2122 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2124 = _T_2122 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2125 = _T_2122 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2126 = regs_10_10 + regs_10_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2146 = {{1'd0}, regs_10_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2127 = _T_2126 + _GEN_2146; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2147 = {{2'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2128 = _T_2127 + _GEN_2147; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2148 = {{3'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2129 = _T_2128 + _GEN_2148; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2149 = {{4'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2130 = _T_2129 + _GEN_2149; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2150 = {{5'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2131 = _T_2130 + _GEN_2150; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2151 = {{6'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2132 = _T_2131 + _GEN_2151; // @[Conwaylife.scala 31:34]
  wire  _T_2133 = _T_2132 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2134 = _T_2132 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2135 = _T_2132 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2136 = regs_10_11 + regs_10_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2152 = {{1'd0}, regs_10_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2137 = _T_2136 + _GEN_2152; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2153 = {{2'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2138 = _T_2137 + _GEN_2153; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2154 = {{3'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2139 = _T_2138 + _GEN_2154; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2155 = {{4'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2140 = _T_2139 + _GEN_2155; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2156 = {{5'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2141 = _T_2140 + _GEN_2156; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2157 = {{6'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2142 = _T_2141 + _GEN_2157; // @[Conwaylife.scala 31:34]
  wire  _T_2143 = _T_2142 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2144 = _T_2142 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2145 = _T_2142 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2146 = regs_10_12 + regs_10_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2158 = {{1'd0}, regs_10_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2147 = _T_2146 + _GEN_2158; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2159 = {{2'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2148 = _T_2147 + _GEN_2159; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2160 = {{3'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2149 = _T_2148 + _GEN_2160; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2161 = {{4'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2150 = _T_2149 + _GEN_2161; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2162 = {{5'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2151 = _T_2150 + _GEN_2162; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2163 = {{6'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2152 = _T_2151 + _GEN_2163; // @[Conwaylife.scala 31:34]
  wire  _T_2153 = _T_2152 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2154 = _T_2152 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2155 = _T_2152 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2156 = regs_10_13 + regs_10_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2164 = {{1'd0}, regs_10_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2157 = _T_2156 + _GEN_2164; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2165 = {{2'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2158 = _T_2157 + _GEN_2165; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2166 = {{3'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2159 = _T_2158 + _GEN_2166; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2167 = {{4'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2160 = _T_2159 + _GEN_2167; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2168 = {{5'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2161 = _T_2160 + _GEN_2168; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2169 = {{6'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2162 = _T_2161 + _GEN_2169; // @[Conwaylife.scala 31:34]
  wire  _T_2163 = _T_2162 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2164 = _T_2162 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2165 = _T_2162 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2166 = regs_10_14 + regs_10_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2170 = {{1'd0}, regs_10_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2167 = _T_2166 + _GEN_2170; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2171 = {{2'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2168 = _T_2167 + _GEN_2171; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2172 = {{3'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2169 = _T_2168 + _GEN_2172; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2173 = {{4'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2170 = _T_2169 + _GEN_2173; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2174 = {{5'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2171 = _T_2170 + _GEN_2174; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2175 = {{6'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2172 = _T_2171 + _GEN_2175; // @[Conwaylife.scala 31:34]
  wire  _T_2173 = _T_2172 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2174 = _T_2172 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2175 = _T_2172 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2176 = regs_11_15 + regs_11_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2176 = {{1'd0}, regs_11_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2177 = _T_2176 + _GEN_2176; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2177 = {{2'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2178 = _T_2177 + _GEN_2177; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2178 = {{3'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2179 = _T_2178 + _GEN_2178; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2179 = {{4'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2180 = _T_2179 + _GEN_2179; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2180 = {{5'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2181 = _T_2180 + _GEN_2180; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2181 = {{6'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2182 = _T_2181 + _GEN_2181; // @[Conwaylife.scala 31:34]
  wire  _T_2183 = _T_2182 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2184 = _T_2182 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2185 = _T_2182 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2186 = regs_11_0 + regs_11_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2182 = {{1'd0}, regs_11_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2187 = _T_2186 + _GEN_2182; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2183 = {{2'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2188 = _T_2187 + _GEN_2183; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2184 = {{3'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2189 = _T_2188 + _GEN_2184; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2185 = {{4'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2190 = _T_2189 + _GEN_2185; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2186 = {{5'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2191 = _T_2190 + _GEN_2186; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2187 = {{6'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2192 = _T_2191 + _GEN_2187; // @[Conwaylife.scala 31:34]
  wire  _T_2193 = _T_2192 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2194 = _T_2192 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2195 = _T_2192 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2196 = regs_11_1 + regs_11_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2188 = {{1'd0}, regs_11_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2197 = _T_2196 + _GEN_2188; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2189 = {{2'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2198 = _T_2197 + _GEN_2189; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2190 = {{3'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2199 = _T_2198 + _GEN_2190; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2191 = {{4'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2200 = _T_2199 + _GEN_2191; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2192 = {{5'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2201 = _T_2200 + _GEN_2192; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2193 = {{6'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2202 = _T_2201 + _GEN_2193; // @[Conwaylife.scala 31:34]
  wire  _T_2203 = _T_2202 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2204 = _T_2202 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2205 = _T_2202 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2206 = regs_11_2 + regs_11_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2194 = {{1'd0}, regs_11_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2207 = _T_2206 + _GEN_2194; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2195 = {{2'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2208 = _T_2207 + _GEN_2195; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2196 = {{3'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2209 = _T_2208 + _GEN_2196; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2197 = {{4'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2210 = _T_2209 + _GEN_2197; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2198 = {{5'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2211 = _T_2210 + _GEN_2198; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2199 = {{6'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2212 = _T_2211 + _GEN_2199; // @[Conwaylife.scala 31:34]
  wire  _T_2213 = _T_2212 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2214 = _T_2212 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2215 = _T_2212 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2216 = regs_11_3 + regs_11_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2200 = {{1'd0}, regs_11_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2217 = _T_2216 + _GEN_2200; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2201 = {{2'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2218 = _T_2217 + _GEN_2201; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2202 = {{3'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2219 = _T_2218 + _GEN_2202; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2203 = {{4'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2220 = _T_2219 + _GEN_2203; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2204 = {{5'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2221 = _T_2220 + _GEN_2204; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2205 = {{6'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2222 = _T_2221 + _GEN_2205; // @[Conwaylife.scala 31:34]
  wire  _T_2223 = _T_2222 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2224 = _T_2222 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2225 = _T_2222 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2226 = regs_11_4 + regs_11_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2206 = {{1'd0}, regs_11_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2227 = _T_2226 + _GEN_2206; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2207 = {{2'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2228 = _T_2227 + _GEN_2207; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2208 = {{3'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2229 = _T_2228 + _GEN_2208; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2209 = {{4'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2230 = _T_2229 + _GEN_2209; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2210 = {{5'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2231 = _T_2230 + _GEN_2210; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2211 = {{6'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2232 = _T_2231 + _GEN_2211; // @[Conwaylife.scala 31:34]
  wire  _T_2233 = _T_2232 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2234 = _T_2232 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2235 = _T_2232 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2236 = regs_11_5 + regs_11_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2212 = {{1'd0}, regs_11_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2237 = _T_2236 + _GEN_2212; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2213 = {{2'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2238 = _T_2237 + _GEN_2213; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2214 = {{3'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2239 = _T_2238 + _GEN_2214; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2215 = {{4'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2240 = _T_2239 + _GEN_2215; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2216 = {{5'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2241 = _T_2240 + _GEN_2216; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2217 = {{6'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2242 = _T_2241 + _GEN_2217; // @[Conwaylife.scala 31:34]
  wire  _T_2243 = _T_2242 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2244 = _T_2242 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2245 = _T_2242 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2246 = regs_11_6 + regs_11_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2218 = {{1'd0}, regs_11_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2247 = _T_2246 + _GEN_2218; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2219 = {{2'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2248 = _T_2247 + _GEN_2219; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2220 = {{3'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2249 = _T_2248 + _GEN_2220; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2221 = {{4'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2250 = _T_2249 + _GEN_2221; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2222 = {{5'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2251 = _T_2250 + _GEN_2222; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2223 = {{6'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2252 = _T_2251 + _GEN_2223; // @[Conwaylife.scala 31:34]
  wire  _T_2253 = _T_2252 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2254 = _T_2252 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2255 = _T_2252 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2256 = regs_11_7 + regs_11_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2224 = {{1'd0}, regs_11_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2257 = _T_2256 + _GEN_2224; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2225 = {{2'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2258 = _T_2257 + _GEN_2225; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2226 = {{3'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2259 = _T_2258 + _GEN_2226; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2227 = {{4'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2260 = _T_2259 + _GEN_2227; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2228 = {{5'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2261 = _T_2260 + _GEN_2228; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2229 = {{6'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2262 = _T_2261 + _GEN_2229; // @[Conwaylife.scala 31:34]
  wire  _T_2263 = _T_2262 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2264 = _T_2262 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2265 = _T_2262 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2266 = regs_11_8 + regs_11_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2230 = {{1'd0}, regs_11_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2267 = _T_2266 + _GEN_2230; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2231 = {{2'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2268 = _T_2267 + _GEN_2231; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2232 = {{3'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2269 = _T_2268 + _GEN_2232; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2233 = {{4'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2270 = _T_2269 + _GEN_2233; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2234 = {{5'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2271 = _T_2270 + _GEN_2234; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2235 = {{6'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2272 = _T_2271 + _GEN_2235; // @[Conwaylife.scala 31:34]
  wire  _T_2273 = _T_2272 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2274 = _T_2272 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2275 = _T_2272 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2276 = regs_11_9 + regs_11_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2236 = {{1'd0}, regs_11_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2277 = _T_2276 + _GEN_2236; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2237 = {{2'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2278 = _T_2277 + _GEN_2237; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2238 = {{3'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2279 = _T_2278 + _GEN_2238; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2239 = {{4'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2280 = _T_2279 + _GEN_2239; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2240 = {{5'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2281 = _T_2280 + _GEN_2240; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2241 = {{6'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2282 = _T_2281 + _GEN_2241; // @[Conwaylife.scala 31:34]
  wire  _T_2283 = _T_2282 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2284 = _T_2282 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2285 = _T_2282 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2286 = regs_11_10 + regs_11_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2242 = {{1'd0}, regs_11_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2287 = _T_2286 + _GEN_2242; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2243 = {{2'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2288 = _T_2287 + _GEN_2243; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2244 = {{3'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2289 = _T_2288 + _GEN_2244; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2245 = {{4'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2290 = _T_2289 + _GEN_2245; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2246 = {{5'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2291 = _T_2290 + _GEN_2246; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2247 = {{6'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2292 = _T_2291 + _GEN_2247; // @[Conwaylife.scala 31:34]
  wire  _T_2293 = _T_2292 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2294 = _T_2292 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2295 = _T_2292 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2296 = regs_11_11 + regs_11_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2248 = {{1'd0}, regs_11_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2297 = _T_2296 + _GEN_2248; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2249 = {{2'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2298 = _T_2297 + _GEN_2249; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2250 = {{3'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2299 = _T_2298 + _GEN_2250; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2251 = {{4'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2300 = _T_2299 + _GEN_2251; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2252 = {{5'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2301 = _T_2300 + _GEN_2252; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2253 = {{6'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2302 = _T_2301 + _GEN_2253; // @[Conwaylife.scala 31:34]
  wire  _T_2303 = _T_2302 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2304 = _T_2302 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2305 = _T_2302 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2306 = regs_11_12 + regs_11_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2254 = {{1'd0}, regs_11_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2307 = _T_2306 + _GEN_2254; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2255 = {{2'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2308 = _T_2307 + _GEN_2255; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2256 = {{3'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2309 = _T_2308 + _GEN_2256; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2257 = {{4'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2310 = _T_2309 + _GEN_2257; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2258 = {{5'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2311 = _T_2310 + _GEN_2258; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2259 = {{6'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2312 = _T_2311 + _GEN_2259; // @[Conwaylife.scala 31:34]
  wire  _T_2313 = _T_2312 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2314 = _T_2312 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2315 = _T_2312 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2316 = regs_11_13 + regs_11_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2260 = {{1'd0}, regs_11_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2317 = _T_2316 + _GEN_2260; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2261 = {{2'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2318 = _T_2317 + _GEN_2261; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2262 = {{3'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2319 = _T_2318 + _GEN_2262; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2263 = {{4'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2320 = _T_2319 + _GEN_2263; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2264 = {{5'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2321 = _T_2320 + _GEN_2264; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2265 = {{6'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2322 = _T_2321 + _GEN_2265; // @[Conwaylife.scala 31:34]
  wire  _T_2323 = _T_2322 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2324 = _T_2322 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2325 = _T_2322 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2326 = regs_11_14 + regs_11_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2266 = {{1'd0}, regs_11_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2327 = _T_2326 + _GEN_2266; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2267 = {{2'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2328 = _T_2327 + _GEN_2267; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2268 = {{3'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2329 = _T_2328 + _GEN_2268; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2269 = {{4'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2330 = _T_2329 + _GEN_2269; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2270 = {{5'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2331 = _T_2330 + _GEN_2270; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2271 = {{6'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2332 = _T_2331 + _GEN_2271; // @[Conwaylife.scala 31:34]
  wire  _T_2333 = _T_2332 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2334 = _T_2332 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2335 = _T_2332 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2336 = regs_12_15 + regs_12_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2272 = {{1'd0}, regs_12_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2337 = _T_2336 + _GEN_2272; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2273 = {{2'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2338 = _T_2337 + _GEN_2273; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2274 = {{3'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2339 = _T_2338 + _GEN_2274; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2275 = {{4'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2340 = _T_2339 + _GEN_2275; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2276 = {{5'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2341 = _T_2340 + _GEN_2276; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2277 = {{6'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2342 = _T_2341 + _GEN_2277; // @[Conwaylife.scala 31:34]
  wire  _T_2343 = _T_2342 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2344 = _T_2342 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2345 = _T_2342 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2346 = regs_12_0 + regs_12_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2278 = {{1'd0}, regs_12_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2347 = _T_2346 + _GEN_2278; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2279 = {{2'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2348 = _T_2347 + _GEN_2279; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2280 = {{3'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2349 = _T_2348 + _GEN_2280; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2281 = {{4'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2350 = _T_2349 + _GEN_2281; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2282 = {{5'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2351 = _T_2350 + _GEN_2282; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2283 = {{6'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2352 = _T_2351 + _GEN_2283; // @[Conwaylife.scala 31:34]
  wire  _T_2353 = _T_2352 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2354 = _T_2352 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2355 = _T_2352 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2356 = regs_12_1 + regs_12_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2284 = {{1'd0}, regs_12_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2357 = _T_2356 + _GEN_2284; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2285 = {{2'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2358 = _T_2357 + _GEN_2285; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2286 = {{3'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2359 = _T_2358 + _GEN_2286; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2287 = {{4'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2360 = _T_2359 + _GEN_2287; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2288 = {{5'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2361 = _T_2360 + _GEN_2288; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2289 = {{6'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2362 = _T_2361 + _GEN_2289; // @[Conwaylife.scala 31:34]
  wire  _T_2363 = _T_2362 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2364 = _T_2362 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2365 = _T_2362 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2366 = regs_12_2 + regs_12_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2290 = {{1'd0}, regs_12_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2367 = _T_2366 + _GEN_2290; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2291 = {{2'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2368 = _T_2367 + _GEN_2291; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2292 = {{3'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2369 = _T_2368 + _GEN_2292; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2293 = {{4'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2370 = _T_2369 + _GEN_2293; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2294 = {{5'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2371 = _T_2370 + _GEN_2294; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2295 = {{6'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2372 = _T_2371 + _GEN_2295; // @[Conwaylife.scala 31:34]
  wire  _T_2373 = _T_2372 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2374 = _T_2372 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2375 = _T_2372 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2376 = regs_12_3 + regs_12_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2296 = {{1'd0}, regs_12_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2377 = _T_2376 + _GEN_2296; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2297 = {{2'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2378 = _T_2377 + _GEN_2297; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2298 = {{3'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2379 = _T_2378 + _GEN_2298; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2299 = {{4'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2380 = _T_2379 + _GEN_2299; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2300 = {{5'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2381 = _T_2380 + _GEN_2300; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2301 = {{6'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2382 = _T_2381 + _GEN_2301; // @[Conwaylife.scala 31:34]
  wire  _T_2383 = _T_2382 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2384 = _T_2382 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2385 = _T_2382 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2386 = regs_12_4 + regs_12_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2302 = {{1'd0}, regs_12_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2387 = _T_2386 + _GEN_2302; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2303 = {{2'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2388 = _T_2387 + _GEN_2303; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2304 = {{3'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2389 = _T_2388 + _GEN_2304; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2305 = {{4'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2390 = _T_2389 + _GEN_2305; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2306 = {{5'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2391 = _T_2390 + _GEN_2306; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2307 = {{6'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2392 = _T_2391 + _GEN_2307; // @[Conwaylife.scala 31:34]
  wire  _T_2393 = _T_2392 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2394 = _T_2392 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2395 = _T_2392 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2396 = regs_12_5 + regs_12_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2308 = {{1'd0}, regs_12_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2397 = _T_2396 + _GEN_2308; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2309 = {{2'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2398 = _T_2397 + _GEN_2309; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2310 = {{3'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2399 = _T_2398 + _GEN_2310; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2311 = {{4'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2400 = _T_2399 + _GEN_2311; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2312 = {{5'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2401 = _T_2400 + _GEN_2312; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2313 = {{6'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2402 = _T_2401 + _GEN_2313; // @[Conwaylife.scala 31:34]
  wire  _T_2403 = _T_2402 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2404 = _T_2402 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2405 = _T_2402 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2406 = regs_12_6 + regs_12_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2314 = {{1'd0}, regs_12_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2407 = _T_2406 + _GEN_2314; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2315 = {{2'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2408 = _T_2407 + _GEN_2315; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2316 = {{3'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2409 = _T_2408 + _GEN_2316; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2317 = {{4'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2410 = _T_2409 + _GEN_2317; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2318 = {{5'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2411 = _T_2410 + _GEN_2318; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2319 = {{6'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2412 = _T_2411 + _GEN_2319; // @[Conwaylife.scala 31:34]
  wire  _T_2413 = _T_2412 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2414 = _T_2412 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2415 = _T_2412 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2416 = regs_12_7 + regs_12_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2320 = {{1'd0}, regs_12_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2417 = _T_2416 + _GEN_2320; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2321 = {{2'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2418 = _T_2417 + _GEN_2321; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2322 = {{3'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2419 = _T_2418 + _GEN_2322; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2323 = {{4'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2420 = _T_2419 + _GEN_2323; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2324 = {{5'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2421 = _T_2420 + _GEN_2324; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2325 = {{6'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2422 = _T_2421 + _GEN_2325; // @[Conwaylife.scala 31:34]
  wire  _T_2423 = _T_2422 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2424 = _T_2422 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2425 = _T_2422 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2426 = regs_12_8 + regs_12_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2326 = {{1'd0}, regs_12_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2427 = _T_2426 + _GEN_2326; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2327 = {{2'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2428 = _T_2427 + _GEN_2327; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2328 = {{3'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2429 = _T_2428 + _GEN_2328; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2329 = {{4'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2430 = _T_2429 + _GEN_2329; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2330 = {{5'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2431 = _T_2430 + _GEN_2330; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2331 = {{6'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2432 = _T_2431 + _GEN_2331; // @[Conwaylife.scala 31:34]
  wire  _T_2433 = _T_2432 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2434 = _T_2432 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2435 = _T_2432 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2436 = regs_12_9 + regs_12_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2332 = {{1'd0}, regs_12_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2437 = _T_2436 + _GEN_2332; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2333 = {{2'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2438 = _T_2437 + _GEN_2333; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2334 = {{3'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2439 = _T_2438 + _GEN_2334; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2335 = {{4'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2440 = _T_2439 + _GEN_2335; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2336 = {{5'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2441 = _T_2440 + _GEN_2336; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2337 = {{6'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2442 = _T_2441 + _GEN_2337; // @[Conwaylife.scala 31:34]
  wire  _T_2443 = _T_2442 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2444 = _T_2442 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2445 = _T_2442 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2446 = regs_12_10 + regs_12_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2338 = {{1'd0}, regs_12_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2447 = _T_2446 + _GEN_2338; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2339 = {{2'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2448 = _T_2447 + _GEN_2339; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2340 = {{3'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2449 = _T_2448 + _GEN_2340; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2341 = {{4'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2450 = _T_2449 + _GEN_2341; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2342 = {{5'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2451 = _T_2450 + _GEN_2342; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2343 = {{6'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2452 = _T_2451 + _GEN_2343; // @[Conwaylife.scala 31:34]
  wire  _T_2453 = _T_2452 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2454 = _T_2452 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2455 = _T_2452 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2456 = regs_12_11 + regs_12_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2344 = {{1'd0}, regs_12_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2457 = _T_2456 + _GEN_2344; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2345 = {{2'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2458 = _T_2457 + _GEN_2345; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2346 = {{3'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2459 = _T_2458 + _GEN_2346; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2347 = {{4'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2460 = _T_2459 + _GEN_2347; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2348 = {{5'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2461 = _T_2460 + _GEN_2348; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2349 = {{6'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2462 = _T_2461 + _GEN_2349; // @[Conwaylife.scala 31:34]
  wire  _T_2463 = _T_2462 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2464 = _T_2462 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2465 = _T_2462 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2466 = regs_12_12 + regs_12_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2350 = {{1'd0}, regs_12_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2467 = _T_2466 + _GEN_2350; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2351 = {{2'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2468 = _T_2467 + _GEN_2351; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2352 = {{3'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2469 = _T_2468 + _GEN_2352; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2353 = {{4'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2470 = _T_2469 + _GEN_2353; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2354 = {{5'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2471 = _T_2470 + _GEN_2354; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2355 = {{6'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2472 = _T_2471 + _GEN_2355; // @[Conwaylife.scala 31:34]
  wire  _T_2473 = _T_2472 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2474 = _T_2472 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2475 = _T_2472 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2476 = regs_12_13 + regs_12_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2356 = {{1'd0}, regs_12_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2477 = _T_2476 + _GEN_2356; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2357 = {{2'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2478 = _T_2477 + _GEN_2357; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2358 = {{3'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2479 = _T_2478 + _GEN_2358; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2359 = {{4'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2480 = _T_2479 + _GEN_2359; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2360 = {{5'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2481 = _T_2480 + _GEN_2360; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2361 = {{6'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2482 = _T_2481 + _GEN_2361; // @[Conwaylife.scala 31:34]
  wire  _T_2483 = _T_2482 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2484 = _T_2482 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2485 = _T_2482 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2486 = regs_12_14 + regs_12_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2362 = {{1'd0}, regs_12_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2487 = _T_2486 + _GEN_2362; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2363 = {{2'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2488 = _T_2487 + _GEN_2363; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2364 = {{3'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2489 = _T_2488 + _GEN_2364; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2365 = {{4'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2490 = _T_2489 + _GEN_2365; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2366 = {{5'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2491 = _T_2490 + _GEN_2366; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2367 = {{6'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2492 = _T_2491 + _GEN_2367; // @[Conwaylife.scala 31:34]
  wire  _T_2493 = _T_2492 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2494 = _T_2492 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2495 = _T_2492 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2496 = regs_13_15 + regs_13_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2368 = {{1'd0}, regs_13_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2497 = _T_2496 + _GEN_2368; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2369 = {{2'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2498 = _T_2497 + _GEN_2369; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2370 = {{3'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2499 = _T_2498 + _GEN_2370; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2371 = {{4'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2500 = _T_2499 + _GEN_2371; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2372 = {{5'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2501 = _T_2500 + _GEN_2372; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2373 = {{6'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2502 = _T_2501 + _GEN_2373; // @[Conwaylife.scala 31:34]
  wire  _T_2503 = _T_2502 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2504 = _T_2502 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2505 = _T_2502 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2506 = regs_13_0 + regs_13_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2374 = {{1'd0}, regs_13_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2507 = _T_2506 + _GEN_2374; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2375 = {{2'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2508 = _T_2507 + _GEN_2375; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2376 = {{3'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2509 = _T_2508 + _GEN_2376; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2377 = {{4'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2510 = _T_2509 + _GEN_2377; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2378 = {{5'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2511 = _T_2510 + _GEN_2378; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2379 = {{6'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2512 = _T_2511 + _GEN_2379; // @[Conwaylife.scala 31:34]
  wire  _T_2513 = _T_2512 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2514 = _T_2512 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2515 = _T_2512 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2516 = regs_13_1 + regs_13_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2380 = {{1'd0}, regs_13_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2517 = _T_2516 + _GEN_2380; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2381 = {{2'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2518 = _T_2517 + _GEN_2381; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2382 = {{3'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2519 = _T_2518 + _GEN_2382; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2383 = {{4'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2520 = _T_2519 + _GEN_2383; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2384 = {{5'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2521 = _T_2520 + _GEN_2384; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2385 = {{6'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2522 = _T_2521 + _GEN_2385; // @[Conwaylife.scala 31:34]
  wire  _T_2523 = _T_2522 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2524 = _T_2522 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2525 = _T_2522 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2526 = regs_13_2 + regs_13_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2386 = {{1'd0}, regs_13_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2527 = _T_2526 + _GEN_2386; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2387 = {{2'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2528 = _T_2527 + _GEN_2387; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2388 = {{3'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2529 = _T_2528 + _GEN_2388; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2389 = {{4'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2530 = _T_2529 + _GEN_2389; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2390 = {{5'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2531 = _T_2530 + _GEN_2390; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2391 = {{6'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2532 = _T_2531 + _GEN_2391; // @[Conwaylife.scala 31:34]
  wire  _T_2533 = _T_2532 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2534 = _T_2532 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2535 = _T_2532 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2536 = regs_13_3 + regs_13_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2392 = {{1'd0}, regs_13_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2537 = _T_2536 + _GEN_2392; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2393 = {{2'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2538 = _T_2537 + _GEN_2393; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2394 = {{3'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2539 = _T_2538 + _GEN_2394; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2395 = {{4'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2540 = _T_2539 + _GEN_2395; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2396 = {{5'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2541 = _T_2540 + _GEN_2396; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2397 = {{6'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2542 = _T_2541 + _GEN_2397; // @[Conwaylife.scala 31:34]
  wire  _T_2543 = _T_2542 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2544 = _T_2542 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2545 = _T_2542 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2546 = regs_13_4 + regs_13_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2398 = {{1'd0}, regs_13_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2547 = _T_2546 + _GEN_2398; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2399 = {{2'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2548 = _T_2547 + _GEN_2399; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2400 = {{3'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2549 = _T_2548 + _GEN_2400; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2401 = {{4'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2550 = _T_2549 + _GEN_2401; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2402 = {{5'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2551 = _T_2550 + _GEN_2402; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2403 = {{6'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2552 = _T_2551 + _GEN_2403; // @[Conwaylife.scala 31:34]
  wire  _T_2553 = _T_2552 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2554 = _T_2552 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2555 = _T_2552 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2556 = regs_13_5 + regs_13_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2404 = {{1'd0}, regs_13_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2557 = _T_2556 + _GEN_2404; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2405 = {{2'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2558 = _T_2557 + _GEN_2405; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2406 = {{3'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2559 = _T_2558 + _GEN_2406; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2407 = {{4'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2560 = _T_2559 + _GEN_2407; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2408 = {{5'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2561 = _T_2560 + _GEN_2408; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2409 = {{6'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2562 = _T_2561 + _GEN_2409; // @[Conwaylife.scala 31:34]
  wire  _T_2563 = _T_2562 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2564 = _T_2562 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2565 = _T_2562 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2566 = regs_13_6 + regs_13_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2410 = {{1'd0}, regs_13_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2567 = _T_2566 + _GEN_2410; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2411 = {{2'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2568 = _T_2567 + _GEN_2411; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2412 = {{3'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2569 = _T_2568 + _GEN_2412; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2413 = {{4'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2570 = _T_2569 + _GEN_2413; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2414 = {{5'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2571 = _T_2570 + _GEN_2414; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2415 = {{6'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2572 = _T_2571 + _GEN_2415; // @[Conwaylife.scala 31:34]
  wire  _T_2573 = _T_2572 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2574 = _T_2572 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2575 = _T_2572 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2576 = regs_13_7 + regs_13_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2416 = {{1'd0}, regs_13_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2577 = _T_2576 + _GEN_2416; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2417 = {{2'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2578 = _T_2577 + _GEN_2417; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2418 = {{3'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2579 = _T_2578 + _GEN_2418; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2419 = {{4'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2580 = _T_2579 + _GEN_2419; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2420 = {{5'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2581 = _T_2580 + _GEN_2420; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2421 = {{6'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2582 = _T_2581 + _GEN_2421; // @[Conwaylife.scala 31:34]
  wire  _T_2583 = _T_2582 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2584 = _T_2582 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2585 = _T_2582 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2586 = regs_13_8 + regs_13_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2422 = {{1'd0}, regs_13_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2587 = _T_2586 + _GEN_2422; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2423 = {{2'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2588 = _T_2587 + _GEN_2423; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2424 = {{3'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2589 = _T_2588 + _GEN_2424; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2425 = {{4'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2590 = _T_2589 + _GEN_2425; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2426 = {{5'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2591 = _T_2590 + _GEN_2426; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2427 = {{6'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2592 = _T_2591 + _GEN_2427; // @[Conwaylife.scala 31:34]
  wire  _T_2593 = _T_2592 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2594 = _T_2592 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2595 = _T_2592 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2596 = regs_13_9 + regs_13_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2428 = {{1'd0}, regs_13_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2597 = _T_2596 + _GEN_2428; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2429 = {{2'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2598 = _T_2597 + _GEN_2429; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2430 = {{3'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2599 = _T_2598 + _GEN_2430; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2431 = {{4'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2600 = _T_2599 + _GEN_2431; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2432 = {{5'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2601 = _T_2600 + _GEN_2432; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2433 = {{6'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2602 = _T_2601 + _GEN_2433; // @[Conwaylife.scala 31:34]
  wire  _T_2603 = _T_2602 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2604 = _T_2602 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2605 = _T_2602 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2606 = regs_13_10 + regs_13_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2434 = {{1'd0}, regs_13_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2607 = _T_2606 + _GEN_2434; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2435 = {{2'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2608 = _T_2607 + _GEN_2435; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2436 = {{3'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2609 = _T_2608 + _GEN_2436; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2437 = {{4'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2610 = _T_2609 + _GEN_2437; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2438 = {{5'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2611 = _T_2610 + _GEN_2438; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2439 = {{6'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2612 = _T_2611 + _GEN_2439; // @[Conwaylife.scala 31:34]
  wire  _T_2613 = _T_2612 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2614 = _T_2612 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2615 = _T_2612 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2616 = regs_13_11 + regs_13_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2440 = {{1'd0}, regs_13_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2617 = _T_2616 + _GEN_2440; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2441 = {{2'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2618 = _T_2617 + _GEN_2441; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2442 = {{3'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2619 = _T_2618 + _GEN_2442; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2443 = {{4'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2620 = _T_2619 + _GEN_2443; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2444 = {{5'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2621 = _T_2620 + _GEN_2444; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2445 = {{6'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2622 = _T_2621 + _GEN_2445; // @[Conwaylife.scala 31:34]
  wire  _T_2623 = _T_2622 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2624 = _T_2622 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2625 = _T_2622 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2626 = regs_13_12 + regs_13_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2446 = {{1'd0}, regs_13_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2627 = _T_2626 + _GEN_2446; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2447 = {{2'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2628 = _T_2627 + _GEN_2447; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2448 = {{3'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2629 = _T_2628 + _GEN_2448; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2449 = {{4'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2630 = _T_2629 + _GEN_2449; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2450 = {{5'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2631 = _T_2630 + _GEN_2450; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2451 = {{6'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2632 = _T_2631 + _GEN_2451; // @[Conwaylife.scala 31:34]
  wire  _T_2633 = _T_2632 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2634 = _T_2632 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2635 = _T_2632 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2636 = regs_13_13 + regs_13_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2452 = {{1'd0}, regs_13_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2637 = _T_2636 + _GEN_2452; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2453 = {{2'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2638 = _T_2637 + _GEN_2453; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2454 = {{3'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2639 = _T_2638 + _GEN_2454; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2455 = {{4'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2640 = _T_2639 + _GEN_2455; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2456 = {{5'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2641 = _T_2640 + _GEN_2456; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2457 = {{6'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2642 = _T_2641 + _GEN_2457; // @[Conwaylife.scala 31:34]
  wire  _T_2643 = _T_2642 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2644 = _T_2642 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2645 = _T_2642 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2646 = regs_13_14 + regs_13_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2458 = {{1'd0}, regs_13_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2647 = _T_2646 + _GEN_2458; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2459 = {{2'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2648 = _T_2647 + _GEN_2459; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2460 = {{3'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2649 = _T_2648 + _GEN_2460; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2461 = {{4'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2650 = _T_2649 + _GEN_2461; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2462 = {{5'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2651 = _T_2650 + _GEN_2462; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2463 = {{6'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2652 = _T_2651 + _GEN_2463; // @[Conwaylife.scala 31:34]
  wire  _T_2653 = _T_2652 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2654 = _T_2652 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2655 = _T_2652 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2656 = regs_14_15 + regs_14_0; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2464 = {{1'd0}, regs_14_1}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2657 = _T_2656 + _GEN_2464; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2465 = {{2'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2658 = _T_2657 + _GEN_2465; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2466 = {{3'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2659 = _T_2658 + _GEN_2466; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2467 = {{4'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2660 = _T_2659 + _GEN_2467; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2468 = {{5'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2661 = _T_2660 + _GEN_2468; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2469 = {{6'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2662 = _T_2661 + _GEN_2469; // @[Conwaylife.scala 31:34]
  wire  _T_2663 = _T_2662 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2664 = _T_2662 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2665 = _T_2662 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2666 = regs_14_0 + regs_14_1; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2470 = {{1'd0}, regs_14_2}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2667 = _T_2666 + _GEN_2470; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2471 = {{2'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2668 = _T_2667 + _GEN_2471; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2472 = {{3'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2669 = _T_2668 + _GEN_2472; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2473 = {{4'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2670 = _T_2669 + _GEN_2473; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2474 = {{5'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2671 = _T_2670 + _GEN_2474; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2475 = {{6'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2672 = _T_2671 + _GEN_2475; // @[Conwaylife.scala 31:34]
  wire  _T_2673 = _T_2672 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2674 = _T_2672 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2675 = _T_2672 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2676 = regs_14_1 + regs_14_2; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2476 = {{1'd0}, regs_14_3}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2677 = _T_2676 + _GEN_2476; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2477 = {{2'd0}, regs_15_1}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2678 = _T_2677 + _GEN_2477; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2478 = {{3'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2679 = _T_2678 + _GEN_2478; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2479 = {{4'd0}, regs_0_1}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2680 = _T_2679 + _GEN_2479; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2480 = {{5'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2681 = _T_2680 + _GEN_2480; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2481 = {{6'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2682 = _T_2681 + _GEN_2481; // @[Conwaylife.scala 31:34]
  wire  _T_2683 = _T_2682 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2684 = _T_2682 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2685 = _T_2682 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2686 = regs_14_2 + regs_14_3; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2482 = {{1'd0}, regs_14_4}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2687 = _T_2686 + _GEN_2482; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2483 = {{2'd0}, regs_15_2}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2688 = _T_2687 + _GEN_2483; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2484 = {{3'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2689 = _T_2688 + _GEN_2484; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2485 = {{4'd0}, regs_0_2}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2690 = _T_2689 + _GEN_2485; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2486 = {{5'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2691 = _T_2690 + _GEN_2486; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2487 = {{6'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2692 = _T_2691 + _GEN_2487; // @[Conwaylife.scala 31:34]
  wire  _T_2693 = _T_2692 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2694 = _T_2692 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2695 = _T_2692 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2696 = regs_14_3 + regs_14_4; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2488 = {{1'd0}, regs_14_5}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2697 = _T_2696 + _GEN_2488; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2489 = {{2'd0}, regs_15_3}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2698 = _T_2697 + _GEN_2489; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2490 = {{3'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2699 = _T_2698 + _GEN_2490; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2491 = {{4'd0}, regs_0_3}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2700 = _T_2699 + _GEN_2491; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2492 = {{5'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2701 = _T_2700 + _GEN_2492; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2493 = {{6'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2702 = _T_2701 + _GEN_2493; // @[Conwaylife.scala 31:34]
  wire  _T_2703 = _T_2702 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2704 = _T_2702 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2705 = _T_2702 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2706 = regs_14_4 + regs_14_5; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2494 = {{1'd0}, regs_14_6}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2707 = _T_2706 + _GEN_2494; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2495 = {{2'd0}, regs_15_4}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2708 = _T_2707 + _GEN_2495; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2496 = {{3'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2709 = _T_2708 + _GEN_2496; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2497 = {{4'd0}, regs_0_4}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2710 = _T_2709 + _GEN_2497; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2498 = {{5'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2711 = _T_2710 + _GEN_2498; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2499 = {{6'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2712 = _T_2711 + _GEN_2499; // @[Conwaylife.scala 31:34]
  wire  _T_2713 = _T_2712 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2714 = _T_2712 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2715 = _T_2712 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2716 = regs_14_5 + regs_14_6; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2500 = {{1'd0}, regs_14_7}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2717 = _T_2716 + _GEN_2500; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2501 = {{2'd0}, regs_15_5}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2718 = _T_2717 + _GEN_2501; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2502 = {{3'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2719 = _T_2718 + _GEN_2502; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2503 = {{4'd0}, regs_0_5}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2720 = _T_2719 + _GEN_2503; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2504 = {{5'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2721 = _T_2720 + _GEN_2504; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2505 = {{6'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2722 = _T_2721 + _GEN_2505; // @[Conwaylife.scala 31:34]
  wire  _T_2723 = _T_2722 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2724 = _T_2722 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2725 = _T_2722 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2726 = regs_14_6 + regs_14_7; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2506 = {{1'd0}, regs_14_8}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2727 = _T_2726 + _GEN_2506; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2507 = {{2'd0}, regs_15_6}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2728 = _T_2727 + _GEN_2507; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2508 = {{3'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2729 = _T_2728 + _GEN_2508; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2509 = {{4'd0}, regs_0_6}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2730 = _T_2729 + _GEN_2509; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2510 = {{5'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2731 = _T_2730 + _GEN_2510; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2511 = {{6'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2732 = _T_2731 + _GEN_2511; // @[Conwaylife.scala 31:34]
  wire  _T_2733 = _T_2732 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2734 = _T_2732 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2735 = _T_2732 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2736 = regs_14_7 + regs_14_8; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2512 = {{1'd0}, regs_14_9}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2737 = _T_2736 + _GEN_2512; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2513 = {{2'd0}, regs_15_7}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2738 = _T_2737 + _GEN_2513; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2514 = {{3'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2739 = _T_2738 + _GEN_2514; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2515 = {{4'd0}, regs_0_7}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2740 = _T_2739 + _GEN_2515; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2516 = {{5'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2741 = _T_2740 + _GEN_2516; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2517 = {{6'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2742 = _T_2741 + _GEN_2517; // @[Conwaylife.scala 31:34]
  wire  _T_2743 = _T_2742 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2744 = _T_2742 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2745 = _T_2742 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2746 = regs_14_8 + regs_14_9; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2518 = {{1'd0}, regs_14_10}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2747 = _T_2746 + _GEN_2518; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2519 = {{2'd0}, regs_15_8}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2748 = _T_2747 + _GEN_2519; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2520 = {{3'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2749 = _T_2748 + _GEN_2520; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2521 = {{4'd0}, regs_0_8}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2750 = _T_2749 + _GEN_2521; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2522 = {{5'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2751 = _T_2750 + _GEN_2522; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2523 = {{6'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2752 = _T_2751 + _GEN_2523; // @[Conwaylife.scala 31:34]
  wire  _T_2753 = _T_2752 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2754 = _T_2752 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2755 = _T_2752 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2756 = regs_14_9 + regs_14_10; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2524 = {{1'd0}, regs_14_11}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2757 = _T_2756 + _GEN_2524; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2525 = {{2'd0}, regs_15_9}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2758 = _T_2757 + _GEN_2525; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2526 = {{3'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2759 = _T_2758 + _GEN_2526; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2527 = {{4'd0}, regs_0_9}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2760 = _T_2759 + _GEN_2527; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2528 = {{5'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2761 = _T_2760 + _GEN_2528; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2529 = {{6'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2762 = _T_2761 + _GEN_2529; // @[Conwaylife.scala 31:34]
  wire  _T_2763 = _T_2762 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2764 = _T_2762 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2765 = _T_2762 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2766 = regs_14_10 + regs_14_11; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2530 = {{1'd0}, regs_14_12}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2767 = _T_2766 + _GEN_2530; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2531 = {{2'd0}, regs_15_10}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2768 = _T_2767 + _GEN_2531; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2532 = {{3'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2769 = _T_2768 + _GEN_2532; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2533 = {{4'd0}, regs_0_10}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2770 = _T_2769 + _GEN_2533; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2534 = {{5'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2771 = _T_2770 + _GEN_2534; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2535 = {{6'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2772 = _T_2771 + _GEN_2535; // @[Conwaylife.scala 31:34]
  wire  _T_2773 = _T_2772 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2774 = _T_2772 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2775 = _T_2772 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2776 = regs_14_11 + regs_14_12; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2536 = {{1'd0}, regs_14_13}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2777 = _T_2776 + _GEN_2536; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2537 = {{2'd0}, regs_15_11}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2778 = _T_2777 + _GEN_2537; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2538 = {{3'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2779 = _T_2778 + _GEN_2538; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2539 = {{4'd0}, regs_0_11}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2780 = _T_2779 + _GEN_2539; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2540 = {{5'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2781 = _T_2780 + _GEN_2540; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2541 = {{6'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2782 = _T_2781 + _GEN_2541; // @[Conwaylife.scala 31:34]
  wire  _T_2783 = _T_2782 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2784 = _T_2782 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2785 = _T_2782 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2786 = regs_14_12 + regs_14_13; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2542 = {{1'd0}, regs_14_14}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2787 = _T_2786 + _GEN_2542; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2543 = {{2'd0}, regs_15_12}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2788 = _T_2787 + _GEN_2543; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2544 = {{3'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2789 = _T_2788 + _GEN_2544; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2545 = {{4'd0}, regs_0_12}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2790 = _T_2789 + _GEN_2545; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2546 = {{5'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2791 = _T_2790 + _GEN_2546; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2547 = {{6'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2792 = _T_2791 + _GEN_2547; // @[Conwaylife.scala 31:34]
  wire  _T_2793 = _T_2792 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2794 = _T_2792 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2795 = _T_2792 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2796 = regs_14_13 + regs_14_14; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2548 = {{1'd0}, regs_14_15}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2797 = _T_2796 + _GEN_2548; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2549 = {{2'd0}, regs_15_13}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2798 = _T_2797 + _GEN_2549; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2550 = {{3'd0}, regs_15_15}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2799 = _T_2798 + _GEN_2550; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2551 = {{4'd0}, regs_0_13}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2800 = _T_2799 + _GEN_2551; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2552 = {{5'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2801 = _T_2800 + _GEN_2552; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2553 = {{6'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2802 = _T_2801 + _GEN_2553; // @[Conwaylife.scala 31:34]
  wire  _T_2803 = _T_2802 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2804 = _T_2802 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2805 = _T_2802 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [1:0] _T_2806 = regs_14_14 + regs_14_15; // @[Conwaylife.scala 31:34]
  wire [1:0] _GEN_2554 = {{1'd0}, regs_14_0}; // @[Conwaylife.scala 31:34]
  wire [2:0] _T_2807 = _T_2806 + _GEN_2554; // @[Conwaylife.scala 31:34]
  wire [2:0] _GEN_2555 = {{2'd0}, regs_15_14}; // @[Conwaylife.scala 31:34]
  wire [3:0] _T_2808 = _T_2807 + _GEN_2555; // @[Conwaylife.scala 31:34]
  wire [3:0] _GEN_2556 = {{3'd0}, regs_15_0}; // @[Conwaylife.scala 31:34]
  wire [4:0] _T_2809 = _T_2808 + _GEN_2556; // @[Conwaylife.scala 31:34]
  wire [4:0] _GEN_2557 = {{4'd0}, regs_0_14}; // @[Conwaylife.scala 31:34]
  wire [5:0] _T_2810 = _T_2809 + _GEN_2557; // @[Conwaylife.scala 31:34]
  wire [5:0] _GEN_2558 = {{5'd0}, regs_0_15}; // @[Conwaylife.scala 31:34]
  wire [6:0] _T_2811 = _T_2810 + _GEN_2558; // @[Conwaylife.scala 31:34]
  wire [6:0] _GEN_2559 = {{6'd0}, regs_0_0}; // @[Conwaylife.scala 31:34]
  wire [7:0] _T_2812 = _T_2811 + _GEN_2559; // @[Conwaylife.scala 31:34]
  wire  _T_2813 = _T_2812 < 8'h2; // @[Conwaylife.scala 33:14]
  wire  _T_2814 = _T_2812 == 8'h2; // @[Conwaylife.scala 35:20]
  wire  _T_2815 = _T_2812 == 8'h3; // @[Conwaylife.scala 37:20]
  wire [7:0] _T_3078 = {regs_0_7,regs_0_6,regs_0_5,regs_0_4,regs_0_3,regs_0_2,regs_0_1,regs_0_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3086 = {regs_0_15,regs_0_14,regs_0_13,regs_0_12,regs_0_11,regs_0_10,regs_0_9,regs_0_8,_T_3078}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3093 = {regs_1_7,regs_1_6,regs_1_5,regs_1_4,regs_1_3,regs_1_2,regs_1_1,regs_1_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3102 = {regs_1_15,regs_1_14,regs_1_13,regs_1_12,regs_1_11,regs_1_10,regs_1_9,regs_1_8,_T_3093,_T_3086}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3109 = {regs_2_7,regs_2_6,regs_2_5,regs_2_4,regs_2_3,regs_2_2,regs_2_1,regs_2_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3117 = {regs_2_15,regs_2_14,regs_2_13,regs_2_12,regs_2_11,regs_2_10,regs_2_9,regs_2_8,_T_3109}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3124 = {regs_3_7,regs_3_6,regs_3_5,regs_3_4,regs_3_3,regs_3_2,regs_3_1,regs_3_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3133 = {regs_3_15,regs_3_14,regs_3_13,regs_3_12,regs_3_11,regs_3_10,regs_3_9,regs_3_8,_T_3124,_T_3117}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3141 = {regs_4_7,regs_4_6,regs_4_5,regs_4_4,regs_4_3,regs_4_2,regs_4_1,regs_4_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3149 = {regs_4_15,regs_4_14,regs_4_13,regs_4_12,regs_4_11,regs_4_10,regs_4_9,regs_4_8,_T_3141}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3156 = {regs_5_7,regs_5_6,regs_5_5,regs_5_4,regs_5_3,regs_5_2,regs_5_1,regs_5_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3165 = {regs_5_15,regs_5_14,regs_5_13,regs_5_12,regs_5_11,regs_5_10,regs_5_9,regs_5_8,_T_3156,_T_3149}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3172 = {regs_6_7,regs_6_6,regs_6_5,regs_6_4,regs_6_3,regs_6_2,regs_6_1,regs_6_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3180 = {regs_6_15,regs_6_14,regs_6_13,regs_6_12,regs_6_11,regs_6_10,regs_6_9,regs_6_8,_T_3172}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3187 = {regs_7_7,regs_7_6,regs_7_5,regs_7_4,regs_7_3,regs_7_2,regs_7_1,regs_7_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3196 = {regs_7_15,regs_7_14,regs_7_13,regs_7_12,regs_7_11,regs_7_10,regs_7_9,regs_7_8,_T_3187,_T_3180}; // @[Conwaylife.scala 47:17]
  wire [127:0] _T_3198 = {_T_3196,_T_3165,_T_3133,_T_3102}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3205 = {regs_8_7,regs_8_6,regs_8_5,regs_8_4,regs_8_3,regs_8_2,regs_8_1,regs_8_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3213 = {regs_8_15,regs_8_14,regs_8_13,regs_8_12,regs_8_11,regs_8_10,regs_8_9,regs_8_8,_T_3205}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3220 = {regs_9_7,regs_9_6,regs_9_5,regs_9_4,regs_9_3,regs_9_2,regs_9_1,regs_9_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3229 = {regs_9_15,regs_9_14,regs_9_13,regs_9_12,regs_9_11,regs_9_10,regs_9_9,regs_9_8,_T_3220,_T_3213}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3236 = {regs_10_7,regs_10_6,regs_10_5,regs_10_4,regs_10_3,regs_10_2,regs_10_1,regs_10_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3244 = {regs_10_15,regs_10_14,regs_10_13,regs_10_12,regs_10_11,regs_10_10,regs_10_9,regs_10_8,_T_3236}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3251 = {regs_11_7,regs_11_6,regs_11_5,regs_11_4,regs_11_3,regs_11_2,regs_11_1,regs_11_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3260 = {regs_11_15,regs_11_14,regs_11_13,regs_11_12,regs_11_11,regs_11_10,regs_11_9,regs_11_8,_T_3251,_T_3244}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3268 = {regs_12_7,regs_12_6,regs_12_5,regs_12_4,regs_12_3,regs_12_2,regs_12_1,regs_12_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3276 = {regs_12_15,regs_12_14,regs_12_13,regs_12_12,regs_12_11,regs_12_10,regs_12_9,regs_12_8,_T_3268}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3283 = {regs_13_7,regs_13_6,regs_13_5,regs_13_4,regs_13_3,regs_13_2,regs_13_1,regs_13_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3292 = {regs_13_15,regs_13_14,regs_13_13,regs_13_12,regs_13_11,regs_13_10,regs_13_9,regs_13_8,_T_3283,_T_3276}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3299 = {regs_14_7,regs_14_6,regs_14_5,regs_14_4,regs_14_3,regs_14_2,regs_14_1,regs_14_0}; // @[Conwaylife.scala 47:17]
  wire [15:0] _T_3307 = {regs_14_15,regs_14_14,regs_14_13,regs_14_12,regs_14_11,regs_14_10,regs_14_9,regs_14_8,_T_3299}; // @[Conwaylife.scala 47:17]
  wire [7:0] _T_3314 = {regs_15_7,regs_15_6,regs_15_5,regs_15_4,regs_15_3,regs_15_2,regs_15_1,regs_15_0}; // @[Conwaylife.scala 47:17]
  wire [31:0] _T_3323 = {regs_15_15,regs_15_14,regs_15_13,regs_15_12,regs_15_11,regs_15_10,regs_15_9,regs_15_8,_T_3314,_T_3307}; // @[Conwaylife.scala 47:17]
  wire [127:0] _T_3325 = {_T_3323,_T_3292,_T_3260,_T_3229}; // @[Conwaylife.scala 47:17]
  assign io_q = {_T_3325,_T_3198}; // @[Conwaylife.scala 47:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  regs_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  regs_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regs_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  regs_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regs_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  regs_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regs_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  regs_0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  regs_0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  regs_0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  regs_0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  regs_0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regs_0_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  regs_0_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  regs_0_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  regs_1_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  regs_1_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  regs_1_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  regs_1_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  regs_1_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  regs_1_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  regs_1_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  regs_1_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  regs_1_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  regs_1_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  regs_1_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  regs_1_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  regs_1_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  regs_1_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  regs_1_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  regs_1_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  regs_2_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  regs_2_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  regs_2_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  regs_2_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  regs_2_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  regs_2_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  regs_2_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  regs_2_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  regs_2_8 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  regs_2_9 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  regs_2_10 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  regs_2_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  regs_2_12 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  regs_2_13 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  regs_2_14 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  regs_2_15 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  regs_3_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  regs_3_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  regs_3_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  regs_3_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  regs_3_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  regs_3_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  regs_3_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  regs_3_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  regs_3_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  regs_3_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  regs_3_10 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  regs_3_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  regs_3_12 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  regs_3_13 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  regs_3_14 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  regs_3_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  regs_4_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  regs_4_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  regs_4_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  regs_4_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  regs_4_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  regs_4_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  regs_4_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  regs_4_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  regs_4_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  regs_4_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  regs_4_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  regs_4_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  regs_4_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  regs_4_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  regs_4_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  regs_4_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  regs_5_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  regs_5_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  regs_5_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  regs_5_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  regs_5_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  regs_5_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  regs_5_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  regs_5_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  regs_5_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  regs_5_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  regs_5_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  regs_5_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  regs_5_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  regs_5_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  regs_5_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  regs_5_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  regs_6_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  regs_6_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  regs_6_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  regs_6_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  regs_6_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  regs_6_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  regs_6_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  regs_6_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  regs_6_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  regs_6_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  regs_6_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  regs_6_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  regs_6_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  regs_6_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  regs_6_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  regs_6_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  regs_7_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  regs_7_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  regs_7_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  regs_7_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  regs_7_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  regs_7_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  regs_7_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  regs_7_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  regs_7_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  regs_7_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  regs_7_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  regs_7_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  regs_7_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  regs_7_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  regs_7_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  regs_7_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  regs_8_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  regs_8_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  regs_8_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  regs_8_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  regs_8_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  regs_8_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  regs_8_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  regs_8_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  regs_8_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  regs_8_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  regs_8_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  regs_8_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  regs_8_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  regs_8_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  regs_8_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  regs_8_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  regs_9_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  regs_9_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  regs_9_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  regs_9_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  regs_9_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  regs_9_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  regs_9_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  regs_9_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  regs_9_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  regs_9_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  regs_9_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  regs_9_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  regs_9_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  regs_9_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  regs_9_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  regs_9_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  regs_10_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  regs_10_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  regs_10_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  regs_10_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  regs_10_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  regs_10_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  regs_10_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  regs_10_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  regs_10_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  regs_10_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  regs_10_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  regs_10_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  regs_10_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  regs_10_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  regs_10_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  regs_10_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  regs_11_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  regs_11_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  regs_11_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  regs_11_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  regs_11_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  regs_11_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  regs_11_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  regs_11_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  regs_11_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  regs_11_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  regs_11_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  regs_11_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  regs_11_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  regs_11_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  regs_11_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  regs_11_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  regs_12_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  regs_12_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  regs_12_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  regs_12_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  regs_12_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  regs_12_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  regs_12_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  regs_12_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  regs_12_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  regs_12_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  regs_12_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  regs_12_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  regs_12_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  regs_12_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  regs_12_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  regs_12_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  regs_13_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  regs_13_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  regs_13_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  regs_13_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  regs_13_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  regs_13_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  regs_13_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  regs_13_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  regs_13_8 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  regs_13_9 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  regs_13_10 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  regs_13_11 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  regs_13_12 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  regs_13_13 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  regs_13_14 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  regs_13_15 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  regs_14_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  regs_14_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  regs_14_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  regs_14_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  regs_14_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  regs_14_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  regs_14_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  regs_14_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  regs_14_8 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  regs_14_9 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  regs_14_10 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  regs_14_11 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  regs_14_12 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  regs_14_13 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  regs_14_14 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  regs_14_15 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  regs_15_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  regs_15_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  regs_15_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  regs_15_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  regs_15_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  regs_15_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  regs_15_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  regs_15_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  regs_15_8 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  regs_15_9 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  regs_15_10 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  regs_15_11 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  regs_15_12 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  regs_15_13 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  regs_15_14 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  regs_15_15 = _RAND_255[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_load) begin
      regs_0_0 <= io_data[0];
    end else if (_T_263) begin
      regs_0_0 <= 1'h0;
    end else if (!(_T_264)) begin
      regs_0_0 <= _T_265;
    end
    if (io_load) begin
      regs_0_1 <= io_data[1];
    end else if (_T_273) begin
      regs_0_1 <= 1'h0;
    end else if (!(_T_274)) begin
      regs_0_1 <= _T_275;
    end
    if (io_load) begin
      regs_0_2 <= io_data[2];
    end else if (_T_283) begin
      regs_0_2 <= 1'h0;
    end else if (!(_T_284)) begin
      regs_0_2 <= _T_285;
    end
    if (io_load) begin
      regs_0_3 <= io_data[3];
    end else if (_T_293) begin
      regs_0_3 <= 1'h0;
    end else if (!(_T_294)) begin
      regs_0_3 <= _T_295;
    end
    if (io_load) begin
      regs_0_4 <= io_data[4];
    end else if (_T_303) begin
      regs_0_4 <= 1'h0;
    end else if (!(_T_304)) begin
      regs_0_4 <= _T_305;
    end
    if (io_load) begin
      regs_0_5 <= io_data[5];
    end else if (_T_313) begin
      regs_0_5 <= 1'h0;
    end else if (!(_T_314)) begin
      regs_0_5 <= _T_315;
    end
    if (io_load) begin
      regs_0_6 <= io_data[6];
    end else if (_T_323) begin
      regs_0_6 <= 1'h0;
    end else if (!(_T_324)) begin
      regs_0_6 <= _T_325;
    end
    if (io_load) begin
      regs_0_7 <= io_data[7];
    end else if (_T_333) begin
      regs_0_7 <= 1'h0;
    end else if (!(_T_334)) begin
      regs_0_7 <= _T_335;
    end
    if (io_load) begin
      regs_0_8 <= io_data[8];
    end else if (_T_343) begin
      regs_0_8 <= 1'h0;
    end else if (!(_T_344)) begin
      regs_0_8 <= _T_345;
    end
    if (io_load) begin
      regs_0_9 <= io_data[9];
    end else if (_T_353) begin
      regs_0_9 <= 1'h0;
    end else if (!(_T_354)) begin
      regs_0_9 <= _T_355;
    end
    if (io_load) begin
      regs_0_10 <= io_data[10];
    end else if (_T_363) begin
      regs_0_10 <= 1'h0;
    end else if (!(_T_364)) begin
      regs_0_10 <= _T_365;
    end
    if (io_load) begin
      regs_0_11 <= io_data[11];
    end else if (_T_373) begin
      regs_0_11 <= 1'h0;
    end else if (!(_T_374)) begin
      regs_0_11 <= _T_375;
    end
    if (io_load) begin
      regs_0_12 <= io_data[12];
    end else if (_T_383) begin
      regs_0_12 <= 1'h0;
    end else if (!(_T_384)) begin
      regs_0_12 <= _T_385;
    end
    if (io_load) begin
      regs_0_13 <= io_data[13];
    end else if (_T_393) begin
      regs_0_13 <= 1'h0;
    end else if (!(_T_394)) begin
      regs_0_13 <= _T_395;
    end
    if (io_load) begin
      regs_0_14 <= io_data[14];
    end else if (_T_403) begin
      regs_0_14 <= 1'h0;
    end else if (!(_T_404)) begin
      regs_0_14 <= _T_405;
    end
    if (io_load) begin
      regs_0_15 <= io_data[15];
    end else if (_T_413) begin
      regs_0_15 <= 1'h0;
    end else if (!(_T_414)) begin
      regs_0_15 <= _T_415;
    end
    if (io_load) begin
      regs_1_0 <= io_data[16];
    end else if (_T_423) begin
      regs_1_0 <= 1'h0;
    end else if (!(_T_424)) begin
      regs_1_0 <= _T_425;
    end
    if (io_load) begin
      regs_1_1 <= io_data[17];
    end else if (_T_433) begin
      regs_1_1 <= 1'h0;
    end else if (!(_T_434)) begin
      regs_1_1 <= _T_435;
    end
    if (io_load) begin
      regs_1_2 <= io_data[18];
    end else if (_T_443) begin
      regs_1_2 <= 1'h0;
    end else if (!(_T_444)) begin
      regs_1_2 <= _T_445;
    end
    if (io_load) begin
      regs_1_3 <= io_data[19];
    end else if (_T_453) begin
      regs_1_3 <= 1'h0;
    end else if (!(_T_454)) begin
      regs_1_3 <= _T_455;
    end
    if (io_load) begin
      regs_1_4 <= io_data[20];
    end else if (_T_463) begin
      regs_1_4 <= 1'h0;
    end else if (!(_T_464)) begin
      regs_1_4 <= _T_465;
    end
    if (io_load) begin
      regs_1_5 <= io_data[21];
    end else if (_T_473) begin
      regs_1_5 <= 1'h0;
    end else if (!(_T_474)) begin
      regs_1_5 <= _T_475;
    end
    if (io_load) begin
      regs_1_6 <= io_data[22];
    end else if (_T_483) begin
      regs_1_6 <= 1'h0;
    end else if (!(_T_484)) begin
      regs_1_6 <= _T_485;
    end
    if (io_load) begin
      regs_1_7 <= io_data[23];
    end else if (_T_493) begin
      regs_1_7 <= 1'h0;
    end else if (!(_T_494)) begin
      regs_1_7 <= _T_495;
    end
    if (io_load) begin
      regs_1_8 <= io_data[24];
    end else if (_T_503) begin
      regs_1_8 <= 1'h0;
    end else if (!(_T_504)) begin
      regs_1_8 <= _T_505;
    end
    if (io_load) begin
      regs_1_9 <= io_data[25];
    end else if (_T_513) begin
      regs_1_9 <= 1'h0;
    end else if (!(_T_514)) begin
      regs_1_9 <= _T_515;
    end
    if (io_load) begin
      regs_1_10 <= io_data[26];
    end else if (_T_523) begin
      regs_1_10 <= 1'h0;
    end else if (!(_T_524)) begin
      regs_1_10 <= _T_525;
    end
    if (io_load) begin
      regs_1_11 <= io_data[27];
    end else if (_T_533) begin
      regs_1_11 <= 1'h0;
    end else if (!(_T_534)) begin
      regs_1_11 <= _T_535;
    end
    if (io_load) begin
      regs_1_12 <= io_data[28];
    end else if (_T_543) begin
      regs_1_12 <= 1'h0;
    end else if (!(_T_544)) begin
      regs_1_12 <= _T_545;
    end
    if (io_load) begin
      regs_1_13 <= io_data[29];
    end else if (_T_553) begin
      regs_1_13 <= 1'h0;
    end else if (!(_T_554)) begin
      regs_1_13 <= _T_555;
    end
    if (io_load) begin
      regs_1_14 <= io_data[30];
    end else if (_T_563) begin
      regs_1_14 <= 1'h0;
    end else if (!(_T_564)) begin
      regs_1_14 <= _T_565;
    end
    if (io_load) begin
      regs_1_15 <= io_data[31];
    end else if (_T_573) begin
      regs_1_15 <= 1'h0;
    end else if (!(_T_574)) begin
      regs_1_15 <= _T_575;
    end
    if (io_load) begin
      regs_2_0 <= io_data[32];
    end else if (_T_583) begin
      regs_2_0 <= 1'h0;
    end else if (!(_T_584)) begin
      regs_2_0 <= _T_585;
    end
    if (io_load) begin
      regs_2_1 <= io_data[33];
    end else if (_T_593) begin
      regs_2_1 <= 1'h0;
    end else if (!(_T_594)) begin
      regs_2_1 <= _T_595;
    end
    if (io_load) begin
      regs_2_2 <= io_data[34];
    end else if (_T_603) begin
      regs_2_2 <= 1'h0;
    end else if (!(_T_604)) begin
      regs_2_2 <= _T_605;
    end
    if (io_load) begin
      regs_2_3 <= io_data[35];
    end else if (_T_613) begin
      regs_2_3 <= 1'h0;
    end else if (!(_T_614)) begin
      regs_2_3 <= _T_615;
    end
    if (io_load) begin
      regs_2_4 <= io_data[36];
    end else if (_T_623) begin
      regs_2_4 <= 1'h0;
    end else if (!(_T_624)) begin
      regs_2_4 <= _T_625;
    end
    if (io_load) begin
      regs_2_5 <= io_data[37];
    end else if (_T_633) begin
      regs_2_5 <= 1'h0;
    end else if (!(_T_634)) begin
      regs_2_5 <= _T_635;
    end
    if (io_load) begin
      regs_2_6 <= io_data[38];
    end else if (_T_643) begin
      regs_2_6 <= 1'h0;
    end else if (!(_T_644)) begin
      regs_2_6 <= _T_645;
    end
    if (io_load) begin
      regs_2_7 <= io_data[39];
    end else if (_T_653) begin
      regs_2_7 <= 1'h0;
    end else if (!(_T_654)) begin
      regs_2_7 <= _T_655;
    end
    if (io_load) begin
      regs_2_8 <= io_data[40];
    end else if (_T_663) begin
      regs_2_8 <= 1'h0;
    end else if (!(_T_664)) begin
      regs_2_8 <= _T_665;
    end
    if (io_load) begin
      regs_2_9 <= io_data[41];
    end else if (_T_673) begin
      regs_2_9 <= 1'h0;
    end else if (!(_T_674)) begin
      regs_2_9 <= _T_675;
    end
    if (io_load) begin
      regs_2_10 <= io_data[42];
    end else if (_T_683) begin
      regs_2_10 <= 1'h0;
    end else if (!(_T_684)) begin
      regs_2_10 <= _T_685;
    end
    if (io_load) begin
      regs_2_11 <= io_data[43];
    end else if (_T_693) begin
      regs_2_11 <= 1'h0;
    end else if (!(_T_694)) begin
      regs_2_11 <= _T_695;
    end
    if (io_load) begin
      regs_2_12 <= io_data[44];
    end else if (_T_703) begin
      regs_2_12 <= 1'h0;
    end else if (!(_T_704)) begin
      regs_2_12 <= _T_705;
    end
    if (io_load) begin
      regs_2_13 <= io_data[45];
    end else if (_T_713) begin
      regs_2_13 <= 1'h0;
    end else if (!(_T_714)) begin
      regs_2_13 <= _T_715;
    end
    if (io_load) begin
      regs_2_14 <= io_data[46];
    end else if (_T_723) begin
      regs_2_14 <= 1'h0;
    end else if (!(_T_724)) begin
      regs_2_14 <= _T_725;
    end
    if (io_load) begin
      regs_2_15 <= io_data[47];
    end else if (_T_733) begin
      regs_2_15 <= 1'h0;
    end else if (!(_T_734)) begin
      regs_2_15 <= _T_735;
    end
    if (io_load) begin
      regs_3_0 <= io_data[48];
    end else if (_T_743) begin
      regs_3_0 <= 1'h0;
    end else if (!(_T_744)) begin
      regs_3_0 <= _T_745;
    end
    if (io_load) begin
      regs_3_1 <= io_data[49];
    end else if (_T_753) begin
      regs_3_1 <= 1'h0;
    end else if (!(_T_754)) begin
      regs_3_1 <= _T_755;
    end
    if (io_load) begin
      regs_3_2 <= io_data[50];
    end else if (_T_763) begin
      regs_3_2 <= 1'h0;
    end else if (!(_T_764)) begin
      regs_3_2 <= _T_765;
    end
    if (io_load) begin
      regs_3_3 <= io_data[51];
    end else if (_T_773) begin
      regs_3_3 <= 1'h0;
    end else if (!(_T_774)) begin
      regs_3_3 <= _T_775;
    end
    if (io_load) begin
      regs_3_4 <= io_data[52];
    end else if (_T_783) begin
      regs_3_4 <= 1'h0;
    end else if (!(_T_784)) begin
      regs_3_4 <= _T_785;
    end
    if (io_load) begin
      regs_3_5 <= io_data[53];
    end else if (_T_793) begin
      regs_3_5 <= 1'h0;
    end else if (!(_T_794)) begin
      regs_3_5 <= _T_795;
    end
    if (io_load) begin
      regs_3_6 <= io_data[54];
    end else if (_T_803) begin
      regs_3_6 <= 1'h0;
    end else if (!(_T_804)) begin
      regs_3_6 <= _T_805;
    end
    if (io_load) begin
      regs_3_7 <= io_data[55];
    end else if (_T_813) begin
      regs_3_7 <= 1'h0;
    end else if (!(_T_814)) begin
      regs_3_7 <= _T_815;
    end
    if (io_load) begin
      regs_3_8 <= io_data[56];
    end else if (_T_823) begin
      regs_3_8 <= 1'h0;
    end else if (!(_T_824)) begin
      regs_3_8 <= _T_825;
    end
    if (io_load) begin
      regs_3_9 <= io_data[57];
    end else if (_T_833) begin
      regs_3_9 <= 1'h0;
    end else if (!(_T_834)) begin
      regs_3_9 <= _T_835;
    end
    if (io_load) begin
      regs_3_10 <= io_data[58];
    end else if (_T_843) begin
      regs_3_10 <= 1'h0;
    end else if (!(_T_844)) begin
      regs_3_10 <= _T_845;
    end
    if (io_load) begin
      regs_3_11 <= io_data[59];
    end else if (_T_853) begin
      regs_3_11 <= 1'h0;
    end else if (!(_T_854)) begin
      regs_3_11 <= _T_855;
    end
    if (io_load) begin
      regs_3_12 <= io_data[60];
    end else if (_T_863) begin
      regs_3_12 <= 1'h0;
    end else if (!(_T_864)) begin
      regs_3_12 <= _T_865;
    end
    if (io_load) begin
      regs_3_13 <= io_data[61];
    end else if (_T_873) begin
      regs_3_13 <= 1'h0;
    end else if (!(_T_874)) begin
      regs_3_13 <= _T_875;
    end
    if (io_load) begin
      regs_3_14 <= io_data[62];
    end else if (_T_883) begin
      regs_3_14 <= 1'h0;
    end else if (!(_T_884)) begin
      regs_3_14 <= _T_885;
    end
    if (io_load) begin
      regs_3_15 <= io_data[63];
    end else if (_T_893) begin
      regs_3_15 <= 1'h0;
    end else if (!(_T_894)) begin
      regs_3_15 <= _T_895;
    end
    if (io_load) begin
      regs_4_0 <= io_data[64];
    end else if (_T_903) begin
      regs_4_0 <= 1'h0;
    end else if (!(_T_904)) begin
      regs_4_0 <= _T_905;
    end
    if (io_load) begin
      regs_4_1 <= io_data[65];
    end else if (_T_913) begin
      regs_4_1 <= 1'h0;
    end else if (!(_T_914)) begin
      regs_4_1 <= _T_915;
    end
    if (io_load) begin
      regs_4_2 <= io_data[66];
    end else if (_T_923) begin
      regs_4_2 <= 1'h0;
    end else if (!(_T_924)) begin
      regs_4_2 <= _T_925;
    end
    if (io_load) begin
      regs_4_3 <= io_data[67];
    end else if (_T_933) begin
      regs_4_3 <= 1'h0;
    end else if (!(_T_934)) begin
      regs_4_3 <= _T_935;
    end
    if (io_load) begin
      regs_4_4 <= io_data[68];
    end else if (_T_943) begin
      regs_4_4 <= 1'h0;
    end else if (!(_T_944)) begin
      regs_4_4 <= _T_945;
    end
    if (io_load) begin
      regs_4_5 <= io_data[69];
    end else if (_T_953) begin
      regs_4_5 <= 1'h0;
    end else if (!(_T_954)) begin
      regs_4_5 <= _T_955;
    end
    if (io_load) begin
      regs_4_6 <= io_data[70];
    end else if (_T_963) begin
      regs_4_6 <= 1'h0;
    end else if (!(_T_964)) begin
      regs_4_6 <= _T_965;
    end
    if (io_load) begin
      regs_4_7 <= io_data[71];
    end else if (_T_973) begin
      regs_4_7 <= 1'h0;
    end else if (!(_T_974)) begin
      regs_4_7 <= _T_975;
    end
    if (io_load) begin
      regs_4_8 <= io_data[72];
    end else if (_T_983) begin
      regs_4_8 <= 1'h0;
    end else if (!(_T_984)) begin
      regs_4_8 <= _T_985;
    end
    if (io_load) begin
      regs_4_9 <= io_data[73];
    end else if (_T_993) begin
      regs_4_9 <= 1'h0;
    end else if (!(_T_994)) begin
      regs_4_9 <= _T_995;
    end
    if (io_load) begin
      regs_4_10 <= io_data[74];
    end else if (_T_1003) begin
      regs_4_10 <= 1'h0;
    end else if (!(_T_1004)) begin
      regs_4_10 <= _T_1005;
    end
    if (io_load) begin
      regs_4_11 <= io_data[75];
    end else if (_T_1013) begin
      regs_4_11 <= 1'h0;
    end else if (!(_T_1014)) begin
      regs_4_11 <= _T_1015;
    end
    if (io_load) begin
      regs_4_12 <= io_data[76];
    end else if (_T_1023) begin
      regs_4_12 <= 1'h0;
    end else if (!(_T_1024)) begin
      regs_4_12 <= _T_1025;
    end
    if (io_load) begin
      regs_4_13 <= io_data[77];
    end else if (_T_1033) begin
      regs_4_13 <= 1'h0;
    end else if (!(_T_1034)) begin
      regs_4_13 <= _T_1035;
    end
    if (io_load) begin
      regs_4_14 <= io_data[78];
    end else if (_T_1043) begin
      regs_4_14 <= 1'h0;
    end else if (!(_T_1044)) begin
      regs_4_14 <= _T_1045;
    end
    if (io_load) begin
      regs_4_15 <= io_data[79];
    end else if (_T_1053) begin
      regs_4_15 <= 1'h0;
    end else if (!(_T_1054)) begin
      regs_4_15 <= _T_1055;
    end
    if (io_load) begin
      regs_5_0 <= io_data[80];
    end else if (_T_1063) begin
      regs_5_0 <= 1'h0;
    end else if (!(_T_1064)) begin
      regs_5_0 <= _T_1065;
    end
    if (io_load) begin
      regs_5_1 <= io_data[81];
    end else if (_T_1073) begin
      regs_5_1 <= 1'h0;
    end else if (!(_T_1074)) begin
      regs_5_1 <= _T_1075;
    end
    if (io_load) begin
      regs_5_2 <= io_data[82];
    end else if (_T_1083) begin
      regs_5_2 <= 1'h0;
    end else if (!(_T_1084)) begin
      regs_5_2 <= _T_1085;
    end
    if (io_load) begin
      regs_5_3 <= io_data[83];
    end else if (_T_1093) begin
      regs_5_3 <= 1'h0;
    end else if (!(_T_1094)) begin
      regs_5_3 <= _T_1095;
    end
    if (io_load) begin
      regs_5_4 <= io_data[84];
    end else if (_T_1103) begin
      regs_5_4 <= 1'h0;
    end else if (!(_T_1104)) begin
      regs_5_4 <= _T_1105;
    end
    if (io_load) begin
      regs_5_5 <= io_data[85];
    end else if (_T_1113) begin
      regs_5_5 <= 1'h0;
    end else if (!(_T_1114)) begin
      regs_5_5 <= _T_1115;
    end
    if (io_load) begin
      regs_5_6 <= io_data[86];
    end else if (_T_1123) begin
      regs_5_6 <= 1'h0;
    end else if (!(_T_1124)) begin
      regs_5_6 <= _T_1125;
    end
    if (io_load) begin
      regs_5_7 <= io_data[87];
    end else if (_T_1133) begin
      regs_5_7 <= 1'h0;
    end else if (!(_T_1134)) begin
      regs_5_7 <= _T_1135;
    end
    if (io_load) begin
      regs_5_8 <= io_data[88];
    end else if (_T_1143) begin
      regs_5_8 <= 1'h0;
    end else if (!(_T_1144)) begin
      regs_5_8 <= _T_1145;
    end
    if (io_load) begin
      regs_5_9 <= io_data[89];
    end else if (_T_1153) begin
      regs_5_9 <= 1'h0;
    end else if (!(_T_1154)) begin
      regs_5_9 <= _T_1155;
    end
    if (io_load) begin
      regs_5_10 <= io_data[90];
    end else if (_T_1163) begin
      regs_5_10 <= 1'h0;
    end else if (!(_T_1164)) begin
      regs_5_10 <= _T_1165;
    end
    if (io_load) begin
      regs_5_11 <= io_data[91];
    end else if (_T_1173) begin
      regs_5_11 <= 1'h0;
    end else if (!(_T_1174)) begin
      regs_5_11 <= _T_1175;
    end
    if (io_load) begin
      regs_5_12 <= io_data[92];
    end else if (_T_1183) begin
      regs_5_12 <= 1'h0;
    end else if (!(_T_1184)) begin
      regs_5_12 <= _T_1185;
    end
    if (io_load) begin
      regs_5_13 <= io_data[93];
    end else if (_T_1193) begin
      regs_5_13 <= 1'h0;
    end else if (!(_T_1194)) begin
      regs_5_13 <= _T_1195;
    end
    if (io_load) begin
      regs_5_14 <= io_data[94];
    end else if (_T_1203) begin
      regs_5_14 <= 1'h0;
    end else if (!(_T_1204)) begin
      regs_5_14 <= _T_1205;
    end
    if (io_load) begin
      regs_5_15 <= io_data[95];
    end else if (_T_1213) begin
      regs_5_15 <= 1'h0;
    end else if (!(_T_1214)) begin
      regs_5_15 <= _T_1215;
    end
    if (io_load) begin
      regs_6_0 <= io_data[96];
    end else if (_T_1223) begin
      regs_6_0 <= 1'h0;
    end else if (!(_T_1224)) begin
      regs_6_0 <= _T_1225;
    end
    if (io_load) begin
      regs_6_1 <= io_data[97];
    end else if (_T_1233) begin
      regs_6_1 <= 1'h0;
    end else if (!(_T_1234)) begin
      regs_6_1 <= _T_1235;
    end
    if (io_load) begin
      regs_6_2 <= io_data[98];
    end else if (_T_1243) begin
      regs_6_2 <= 1'h0;
    end else if (!(_T_1244)) begin
      regs_6_2 <= _T_1245;
    end
    if (io_load) begin
      regs_6_3 <= io_data[99];
    end else if (_T_1253) begin
      regs_6_3 <= 1'h0;
    end else if (!(_T_1254)) begin
      regs_6_3 <= _T_1255;
    end
    if (io_load) begin
      regs_6_4 <= io_data[100];
    end else if (_T_1263) begin
      regs_6_4 <= 1'h0;
    end else if (!(_T_1264)) begin
      regs_6_4 <= _T_1265;
    end
    if (io_load) begin
      regs_6_5 <= io_data[101];
    end else if (_T_1273) begin
      regs_6_5 <= 1'h0;
    end else if (!(_T_1274)) begin
      regs_6_5 <= _T_1275;
    end
    if (io_load) begin
      regs_6_6 <= io_data[102];
    end else if (_T_1283) begin
      regs_6_6 <= 1'h0;
    end else if (!(_T_1284)) begin
      regs_6_6 <= _T_1285;
    end
    if (io_load) begin
      regs_6_7 <= io_data[103];
    end else if (_T_1293) begin
      regs_6_7 <= 1'h0;
    end else if (!(_T_1294)) begin
      regs_6_7 <= _T_1295;
    end
    if (io_load) begin
      regs_6_8 <= io_data[104];
    end else if (_T_1303) begin
      regs_6_8 <= 1'h0;
    end else if (!(_T_1304)) begin
      regs_6_8 <= _T_1305;
    end
    if (io_load) begin
      regs_6_9 <= io_data[105];
    end else if (_T_1313) begin
      regs_6_9 <= 1'h0;
    end else if (!(_T_1314)) begin
      regs_6_9 <= _T_1315;
    end
    if (io_load) begin
      regs_6_10 <= io_data[106];
    end else if (_T_1323) begin
      regs_6_10 <= 1'h0;
    end else if (!(_T_1324)) begin
      regs_6_10 <= _T_1325;
    end
    if (io_load) begin
      regs_6_11 <= io_data[107];
    end else if (_T_1333) begin
      regs_6_11 <= 1'h0;
    end else if (!(_T_1334)) begin
      regs_6_11 <= _T_1335;
    end
    if (io_load) begin
      regs_6_12 <= io_data[108];
    end else if (_T_1343) begin
      regs_6_12 <= 1'h0;
    end else if (!(_T_1344)) begin
      regs_6_12 <= _T_1345;
    end
    if (io_load) begin
      regs_6_13 <= io_data[109];
    end else if (_T_1353) begin
      regs_6_13 <= 1'h0;
    end else if (!(_T_1354)) begin
      regs_6_13 <= _T_1355;
    end
    if (io_load) begin
      regs_6_14 <= io_data[110];
    end else if (_T_1363) begin
      regs_6_14 <= 1'h0;
    end else if (!(_T_1364)) begin
      regs_6_14 <= _T_1365;
    end
    if (io_load) begin
      regs_6_15 <= io_data[111];
    end else if (_T_1373) begin
      regs_6_15 <= 1'h0;
    end else if (!(_T_1374)) begin
      regs_6_15 <= _T_1375;
    end
    if (io_load) begin
      regs_7_0 <= io_data[112];
    end else if (_T_1383) begin
      regs_7_0 <= 1'h0;
    end else if (!(_T_1384)) begin
      regs_7_0 <= _T_1385;
    end
    if (io_load) begin
      regs_7_1 <= io_data[113];
    end else if (_T_1393) begin
      regs_7_1 <= 1'h0;
    end else if (!(_T_1394)) begin
      regs_7_1 <= _T_1395;
    end
    if (io_load) begin
      regs_7_2 <= io_data[114];
    end else if (_T_1403) begin
      regs_7_2 <= 1'h0;
    end else if (!(_T_1404)) begin
      regs_7_2 <= _T_1405;
    end
    if (io_load) begin
      regs_7_3 <= io_data[115];
    end else if (_T_1413) begin
      regs_7_3 <= 1'h0;
    end else if (!(_T_1414)) begin
      regs_7_3 <= _T_1415;
    end
    if (io_load) begin
      regs_7_4 <= io_data[116];
    end else if (_T_1423) begin
      regs_7_4 <= 1'h0;
    end else if (!(_T_1424)) begin
      regs_7_4 <= _T_1425;
    end
    if (io_load) begin
      regs_7_5 <= io_data[117];
    end else if (_T_1433) begin
      regs_7_5 <= 1'h0;
    end else if (!(_T_1434)) begin
      regs_7_5 <= _T_1435;
    end
    if (io_load) begin
      regs_7_6 <= io_data[118];
    end else if (_T_1443) begin
      regs_7_6 <= 1'h0;
    end else if (!(_T_1444)) begin
      regs_7_6 <= _T_1445;
    end
    if (io_load) begin
      regs_7_7 <= io_data[119];
    end else if (_T_1453) begin
      regs_7_7 <= 1'h0;
    end else if (!(_T_1454)) begin
      regs_7_7 <= _T_1455;
    end
    if (io_load) begin
      regs_7_8 <= io_data[120];
    end else if (_T_1463) begin
      regs_7_8 <= 1'h0;
    end else if (!(_T_1464)) begin
      regs_7_8 <= _T_1465;
    end
    if (io_load) begin
      regs_7_9 <= io_data[121];
    end else if (_T_1473) begin
      regs_7_9 <= 1'h0;
    end else if (!(_T_1474)) begin
      regs_7_9 <= _T_1475;
    end
    if (io_load) begin
      regs_7_10 <= io_data[122];
    end else if (_T_1483) begin
      regs_7_10 <= 1'h0;
    end else if (!(_T_1484)) begin
      regs_7_10 <= _T_1485;
    end
    if (io_load) begin
      regs_7_11 <= io_data[123];
    end else if (_T_1493) begin
      regs_7_11 <= 1'h0;
    end else if (!(_T_1494)) begin
      regs_7_11 <= _T_1495;
    end
    if (io_load) begin
      regs_7_12 <= io_data[124];
    end else if (_T_1503) begin
      regs_7_12 <= 1'h0;
    end else if (!(_T_1504)) begin
      regs_7_12 <= _T_1505;
    end
    if (io_load) begin
      regs_7_13 <= io_data[125];
    end else if (_T_1513) begin
      regs_7_13 <= 1'h0;
    end else if (!(_T_1514)) begin
      regs_7_13 <= _T_1515;
    end
    if (io_load) begin
      regs_7_14 <= io_data[126];
    end else if (_T_1523) begin
      regs_7_14 <= 1'h0;
    end else if (!(_T_1524)) begin
      regs_7_14 <= _T_1525;
    end
    if (io_load) begin
      regs_7_15 <= io_data[127];
    end else if (_T_1533) begin
      regs_7_15 <= 1'h0;
    end else if (!(_T_1534)) begin
      regs_7_15 <= _T_1535;
    end
    if (io_load) begin
      regs_8_0 <= io_data[128];
    end else if (_T_1543) begin
      regs_8_0 <= 1'h0;
    end else if (!(_T_1544)) begin
      regs_8_0 <= _T_1545;
    end
    if (io_load) begin
      regs_8_1 <= io_data[129];
    end else if (_T_1553) begin
      regs_8_1 <= 1'h0;
    end else if (!(_T_1554)) begin
      regs_8_1 <= _T_1555;
    end
    if (io_load) begin
      regs_8_2 <= io_data[130];
    end else if (_T_1563) begin
      regs_8_2 <= 1'h0;
    end else if (!(_T_1564)) begin
      regs_8_2 <= _T_1565;
    end
    if (io_load) begin
      regs_8_3 <= io_data[131];
    end else if (_T_1573) begin
      regs_8_3 <= 1'h0;
    end else if (!(_T_1574)) begin
      regs_8_3 <= _T_1575;
    end
    if (io_load) begin
      regs_8_4 <= io_data[132];
    end else if (_T_1583) begin
      regs_8_4 <= 1'h0;
    end else if (!(_T_1584)) begin
      regs_8_4 <= _T_1585;
    end
    if (io_load) begin
      regs_8_5 <= io_data[133];
    end else if (_T_1593) begin
      regs_8_5 <= 1'h0;
    end else if (!(_T_1594)) begin
      regs_8_5 <= _T_1595;
    end
    if (io_load) begin
      regs_8_6 <= io_data[134];
    end else if (_T_1603) begin
      regs_8_6 <= 1'h0;
    end else if (!(_T_1604)) begin
      regs_8_6 <= _T_1605;
    end
    if (io_load) begin
      regs_8_7 <= io_data[135];
    end else if (_T_1613) begin
      regs_8_7 <= 1'h0;
    end else if (!(_T_1614)) begin
      regs_8_7 <= _T_1615;
    end
    if (io_load) begin
      regs_8_8 <= io_data[136];
    end else if (_T_1623) begin
      regs_8_8 <= 1'h0;
    end else if (!(_T_1624)) begin
      regs_8_8 <= _T_1625;
    end
    if (io_load) begin
      regs_8_9 <= io_data[137];
    end else if (_T_1633) begin
      regs_8_9 <= 1'h0;
    end else if (!(_T_1634)) begin
      regs_8_9 <= _T_1635;
    end
    if (io_load) begin
      regs_8_10 <= io_data[138];
    end else if (_T_1643) begin
      regs_8_10 <= 1'h0;
    end else if (!(_T_1644)) begin
      regs_8_10 <= _T_1645;
    end
    if (io_load) begin
      regs_8_11 <= io_data[139];
    end else if (_T_1653) begin
      regs_8_11 <= 1'h0;
    end else if (!(_T_1654)) begin
      regs_8_11 <= _T_1655;
    end
    if (io_load) begin
      regs_8_12 <= io_data[140];
    end else if (_T_1663) begin
      regs_8_12 <= 1'h0;
    end else if (!(_T_1664)) begin
      regs_8_12 <= _T_1665;
    end
    if (io_load) begin
      regs_8_13 <= io_data[141];
    end else if (_T_1673) begin
      regs_8_13 <= 1'h0;
    end else if (!(_T_1674)) begin
      regs_8_13 <= _T_1675;
    end
    if (io_load) begin
      regs_8_14 <= io_data[142];
    end else if (_T_1683) begin
      regs_8_14 <= 1'h0;
    end else if (!(_T_1684)) begin
      regs_8_14 <= _T_1685;
    end
    if (io_load) begin
      regs_8_15 <= io_data[143];
    end else if (_T_1693) begin
      regs_8_15 <= 1'h0;
    end else if (!(_T_1694)) begin
      regs_8_15 <= _T_1695;
    end
    if (io_load) begin
      regs_9_0 <= io_data[144];
    end else if (_T_1703) begin
      regs_9_0 <= 1'h0;
    end else if (!(_T_1704)) begin
      regs_9_0 <= _T_1705;
    end
    if (io_load) begin
      regs_9_1 <= io_data[145];
    end else if (_T_1713) begin
      regs_9_1 <= 1'h0;
    end else if (!(_T_1714)) begin
      regs_9_1 <= _T_1715;
    end
    if (io_load) begin
      regs_9_2 <= io_data[146];
    end else if (_T_1723) begin
      regs_9_2 <= 1'h0;
    end else if (!(_T_1724)) begin
      regs_9_2 <= _T_1725;
    end
    if (io_load) begin
      regs_9_3 <= io_data[147];
    end else if (_T_1733) begin
      regs_9_3 <= 1'h0;
    end else if (!(_T_1734)) begin
      regs_9_3 <= _T_1735;
    end
    if (io_load) begin
      regs_9_4 <= io_data[148];
    end else if (_T_1743) begin
      regs_9_4 <= 1'h0;
    end else if (!(_T_1744)) begin
      regs_9_4 <= _T_1745;
    end
    if (io_load) begin
      regs_9_5 <= io_data[149];
    end else if (_T_1753) begin
      regs_9_5 <= 1'h0;
    end else if (!(_T_1754)) begin
      regs_9_5 <= _T_1755;
    end
    if (io_load) begin
      regs_9_6 <= io_data[150];
    end else if (_T_1763) begin
      regs_9_6 <= 1'h0;
    end else if (!(_T_1764)) begin
      regs_9_6 <= _T_1765;
    end
    if (io_load) begin
      regs_9_7 <= io_data[151];
    end else if (_T_1773) begin
      regs_9_7 <= 1'h0;
    end else if (!(_T_1774)) begin
      regs_9_7 <= _T_1775;
    end
    if (io_load) begin
      regs_9_8 <= io_data[152];
    end else if (_T_1783) begin
      regs_9_8 <= 1'h0;
    end else if (!(_T_1784)) begin
      regs_9_8 <= _T_1785;
    end
    if (io_load) begin
      regs_9_9 <= io_data[153];
    end else if (_T_1793) begin
      regs_9_9 <= 1'h0;
    end else if (!(_T_1794)) begin
      regs_9_9 <= _T_1795;
    end
    if (io_load) begin
      regs_9_10 <= io_data[154];
    end else if (_T_1803) begin
      regs_9_10 <= 1'h0;
    end else if (!(_T_1804)) begin
      regs_9_10 <= _T_1805;
    end
    if (io_load) begin
      regs_9_11 <= io_data[155];
    end else if (_T_1813) begin
      regs_9_11 <= 1'h0;
    end else if (!(_T_1814)) begin
      regs_9_11 <= _T_1815;
    end
    if (io_load) begin
      regs_9_12 <= io_data[156];
    end else if (_T_1823) begin
      regs_9_12 <= 1'h0;
    end else if (!(_T_1824)) begin
      regs_9_12 <= _T_1825;
    end
    if (io_load) begin
      regs_9_13 <= io_data[157];
    end else if (_T_1833) begin
      regs_9_13 <= 1'h0;
    end else if (!(_T_1834)) begin
      regs_9_13 <= _T_1835;
    end
    if (io_load) begin
      regs_9_14 <= io_data[158];
    end else if (_T_1843) begin
      regs_9_14 <= 1'h0;
    end else if (!(_T_1844)) begin
      regs_9_14 <= _T_1845;
    end
    if (io_load) begin
      regs_9_15 <= io_data[159];
    end else if (_T_1853) begin
      regs_9_15 <= 1'h0;
    end else if (!(_T_1854)) begin
      regs_9_15 <= _T_1855;
    end
    if (io_load) begin
      regs_10_0 <= io_data[160];
    end else if (_T_1863) begin
      regs_10_0 <= 1'h0;
    end else if (!(_T_1864)) begin
      regs_10_0 <= _T_1865;
    end
    if (io_load) begin
      regs_10_1 <= io_data[161];
    end else if (_T_1873) begin
      regs_10_1 <= 1'h0;
    end else if (!(_T_1874)) begin
      regs_10_1 <= _T_1875;
    end
    if (io_load) begin
      regs_10_2 <= io_data[162];
    end else if (_T_1883) begin
      regs_10_2 <= 1'h0;
    end else if (!(_T_1884)) begin
      regs_10_2 <= _T_1885;
    end
    if (io_load) begin
      regs_10_3 <= io_data[163];
    end else if (_T_1893) begin
      regs_10_3 <= 1'h0;
    end else if (!(_T_1894)) begin
      regs_10_3 <= _T_1895;
    end
    if (io_load) begin
      regs_10_4 <= io_data[164];
    end else if (_T_1903) begin
      regs_10_4 <= 1'h0;
    end else if (!(_T_1904)) begin
      regs_10_4 <= _T_1905;
    end
    if (io_load) begin
      regs_10_5 <= io_data[165];
    end else if (_T_1913) begin
      regs_10_5 <= 1'h0;
    end else if (!(_T_1914)) begin
      regs_10_5 <= _T_1915;
    end
    if (io_load) begin
      regs_10_6 <= io_data[166];
    end else if (_T_1923) begin
      regs_10_6 <= 1'h0;
    end else if (!(_T_1924)) begin
      regs_10_6 <= _T_1925;
    end
    if (io_load) begin
      regs_10_7 <= io_data[167];
    end else if (_T_1933) begin
      regs_10_7 <= 1'h0;
    end else if (!(_T_1934)) begin
      regs_10_7 <= _T_1935;
    end
    if (io_load) begin
      regs_10_8 <= io_data[168];
    end else if (_T_1943) begin
      regs_10_8 <= 1'h0;
    end else if (!(_T_1944)) begin
      regs_10_8 <= _T_1945;
    end
    if (io_load) begin
      regs_10_9 <= io_data[169];
    end else if (_T_1953) begin
      regs_10_9 <= 1'h0;
    end else if (!(_T_1954)) begin
      regs_10_9 <= _T_1955;
    end
    if (io_load) begin
      regs_10_10 <= io_data[170];
    end else if (_T_1963) begin
      regs_10_10 <= 1'h0;
    end else if (!(_T_1964)) begin
      regs_10_10 <= _T_1965;
    end
    if (io_load) begin
      regs_10_11 <= io_data[171];
    end else if (_T_1973) begin
      regs_10_11 <= 1'h0;
    end else if (!(_T_1974)) begin
      regs_10_11 <= _T_1975;
    end
    if (io_load) begin
      regs_10_12 <= io_data[172];
    end else if (_T_1983) begin
      regs_10_12 <= 1'h0;
    end else if (!(_T_1984)) begin
      regs_10_12 <= _T_1985;
    end
    if (io_load) begin
      regs_10_13 <= io_data[173];
    end else if (_T_1993) begin
      regs_10_13 <= 1'h0;
    end else if (!(_T_1994)) begin
      regs_10_13 <= _T_1995;
    end
    if (io_load) begin
      regs_10_14 <= io_data[174];
    end else if (_T_2003) begin
      regs_10_14 <= 1'h0;
    end else if (!(_T_2004)) begin
      regs_10_14 <= _T_2005;
    end
    if (io_load) begin
      regs_10_15 <= io_data[175];
    end else if (_T_2013) begin
      regs_10_15 <= 1'h0;
    end else if (!(_T_2014)) begin
      regs_10_15 <= _T_2015;
    end
    if (io_load) begin
      regs_11_0 <= io_data[176];
    end else if (_T_2023) begin
      regs_11_0 <= 1'h0;
    end else if (!(_T_2024)) begin
      regs_11_0 <= _T_2025;
    end
    if (io_load) begin
      regs_11_1 <= io_data[177];
    end else if (_T_2033) begin
      regs_11_1 <= 1'h0;
    end else if (!(_T_2034)) begin
      regs_11_1 <= _T_2035;
    end
    if (io_load) begin
      regs_11_2 <= io_data[178];
    end else if (_T_2043) begin
      regs_11_2 <= 1'h0;
    end else if (!(_T_2044)) begin
      regs_11_2 <= _T_2045;
    end
    if (io_load) begin
      regs_11_3 <= io_data[179];
    end else if (_T_2053) begin
      regs_11_3 <= 1'h0;
    end else if (!(_T_2054)) begin
      regs_11_3 <= _T_2055;
    end
    if (io_load) begin
      regs_11_4 <= io_data[180];
    end else if (_T_2063) begin
      regs_11_4 <= 1'h0;
    end else if (!(_T_2064)) begin
      regs_11_4 <= _T_2065;
    end
    if (io_load) begin
      regs_11_5 <= io_data[181];
    end else if (_T_2073) begin
      regs_11_5 <= 1'h0;
    end else if (!(_T_2074)) begin
      regs_11_5 <= _T_2075;
    end
    if (io_load) begin
      regs_11_6 <= io_data[182];
    end else if (_T_2083) begin
      regs_11_6 <= 1'h0;
    end else if (!(_T_2084)) begin
      regs_11_6 <= _T_2085;
    end
    if (io_load) begin
      regs_11_7 <= io_data[183];
    end else if (_T_2093) begin
      regs_11_7 <= 1'h0;
    end else if (!(_T_2094)) begin
      regs_11_7 <= _T_2095;
    end
    if (io_load) begin
      regs_11_8 <= io_data[184];
    end else if (_T_2103) begin
      regs_11_8 <= 1'h0;
    end else if (!(_T_2104)) begin
      regs_11_8 <= _T_2105;
    end
    if (io_load) begin
      regs_11_9 <= io_data[185];
    end else if (_T_2113) begin
      regs_11_9 <= 1'h0;
    end else if (!(_T_2114)) begin
      regs_11_9 <= _T_2115;
    end
    if (io_load) begin
      regs_11_10 <= io_data[186];
    end else if (_T_2123) begin
      regs_11_10 <= 1'h0;
    end else if (!(_T_2124)) begin
      regs_11_10 <= _T_2125;
    end
    if (io_load) begin
      regs_11_11 <= io_data[187];
    end else if (_T_2133) begin
      regs_11_11 <= 1'h0;
    end else if (!(_T_2134)) begin
      regs_11_11 <= _T_2135;
    end
    if (io_load) begin
      regs_11_12 <= io_data[188];
    end else if (_T_2143) begin
      regs_11_12 <= 1'h0;
    end else if (!(_T_2144)) begin
      regs_11_12 <= _T_2145;
    end
    if (io_load) begin
      regs_11_13 <= io_data[189];
    end else if (_T_2153) begin
      regs_11_13 <= 1'h0;
    end else if (!(_T_2154)) begin
      regs_11_13 <= _T_2155;
    end
    if (io_load) begin
      regs_11_14 <= io_data[190];
    end else if (_T_2163) begin
      regs_11_14 <= 1'h0;
    end else if (!(_T_2164)) begin
      regs_11_14 <= _T_2165;
    end
    if (io_load) begin
      regs_11_15 <= io_data[191];
    end else if (_T_2173) begin
      regs_11_15 <= 1'h0;
    end else if (!(_T_2174)) begin
      regs_11_15 <= _T_2175;
    end
    if (io_load) begin
      regs_12_0 <= io_data[192];
    end else if (_T_2183) begin
      regs_12_0 <= 1'h0;
    end else if (!(_T_2184)) begin
      regs_12_0 <= _T_2185;
    end
    if (io_load) begin
      regs_12_1 <= io_data[193];
    end else if (_T_2193) begin
      regs_12_1 <= 1'h0;
    end else if (!(_T_2194)) begin
      regs_12_1 <= _T_2195;
    end
    if (io_load) begin
      regs_12_2 <= io_data[194];
    end else if (_T_2203) begin
      regs_12_2 <= 1'h0;
    end else if (!(_T_2204)) begin
      regs_12_2 <= _T_2205;
    end
    if (io_load) begin
      regs_12_3 <= io_data[195];
    end else if (_T_2213) begin
      regs_12_3 <= 1'h0;
    end else if (!(_T_2214)) begin
      regs_12_3 <= _T_2215;
    end
    if (io_load) begin
      regs_12_4 <= io_data[196];
    end else if (_T_2223) begin
      regs_12_4 <= 1'h0;
    end else if (!(_T_2224)) begin
      regs_12_4 <= _T_2225;
    end
    if (io_load) begin
      regs_12_5 <= io_data[197];
    end else if (_T_2233) begin
      regs_12_5 <= 1'h0;
    end else if (!(_T_2234)) begin
      regs_12_5 <= _T_2235;
    end
    if (io_load) begin
      regs_12_6 <= io_data[198];
    end else if (_T_2243) begin
      regs_12_6 <= 1'h0;
    end else if (!(_T_2244)) begin
      regs_12_6 <= _T_2245;
    end
    if (io_load) begin
      regs_12_7 <= io_data[199];
    end else if (_T_2253) begin
      regs_12_7 <= 1'h0;
    end else if (!(_T_2254)) begin
      regs_12_7 <= _T_2255;
    end
    if (io_load) begin
      regs_12_8 <= io_data[200];
    end else if (_T_2263) begin
      regs_12_8 <= 1'h0;
    end else if (!(_T_2264)) begin
      regs_12_8 <= _T_2265;
    end
    if (io_load) begin
      regs_12_9 <= io_data[201];
    end else if (_T_2273) begin
      regs_12_9 <= 1'h0;
    end else if (!(_T_2274)) begin
      regs_12_9 <= _T_2275;
    end
    if (io_load) begin
      regs_12_10 <= io_data[202];
    end else if (_T_2283) begin
      regs_12_10 <= 1'h0;
    end else if (!(_T_2284)) begin
      regs_12_10 <= _T_2285;
    end
    if (io_load) begin
      regs_12_11 <= io_data[203];
    end else if (_T_2293) begin
      regs_12_11 <= 1'h0;
    end else if (!(_T_2294)) begin
      regs_12_11 <= _T_2295;
    end
    if (io_load) begin
      regs_12_12 <= io_data[204];
    end else if (_T_2303) begin
      regs_12_12 <= 1'h0;
    end else if (!(_T_2304)) begin
      regs_12_12 <= _T_2305;
    end
    if (io_load) begin
      regs_12_13 <= io_data[205];
    end else if (_T_2313) begin
      regs_12_13 <= 1'h0;
    end else if (!(_T_2314)) begin
      regs_12_13 <= _T_2315;
    end
    if (io_load) begin
      regs_12_14 <= io_data[206];
    end else if (_T_2323) begin
      regs_12_14 <= 1'h0;
    end else if (!(_T_2324)) begin
      regs_12_14 <= _T_2325;
    end
    if (io_load) begin
      regs_12_15 <= io_data[207];
    end else if (_T_2333) begin
      regs_12_15 <= 1'h0;
    end else if (!(_T_2334)) begin
      regs_12_15 <= _T_2335;
    end
    if (io_load) begin
      regs_13_0 <= io_data[208];
    end else if (_T_2343) begin
      regs_13_0 <= 1'h0;
    end else if (!(_T_2344)) begin
      regs_13_0 <= _T_2345;
    end
    if (io_load) begin
      regs_13_1 <= io_data[209];
    end else if (_T_2353) begin
      regs_13_1 <= 1'h0;
    end else if (!(_T_2354)) begin
      regs_13_1 <= _T_2355;
    end
    if (io_load) begin
      regs_13_2 <= io_data[210];
    end else if (_T_2363) begin
      regs_13_2 <= 1'h0;
    end else if (!(_T_2364)) begin
      regs_13_2 <= _T_2365;
    end
    if (io_load) begin
      regs_13_3 <= io_data[211];
    end else if (_T_2373) begin
      regs_13_3 <= 1'h0;
    end else if (!(_T_2374)) begin
      regs_13_3 <= _T_2375;
    end
    if (io_load) begin
      regs_13_4 <= io_data[212];
    end else if (_T_2383) begin
      regs_13_4 <= 1'h0;
    end else if (!(_T_2384)) begin
      regs_13_4 <= _T_2385;
    end
    if (io_load) begin
      regs_13_5 <= io_data[213];
    end else if (_T_2393) begin
      regs_13_5 <= 1'h0;
    end else if (!(_T_2394)) begin
      regs_13_5 <= _T_2395;
    end
    if (io_load) begin
      regs_13_6 <= io_data[214];
    end else if (_T_2403) begin
      regs_13_6 <= 1'h0;
    end else if (!(_T_2404)) begin
      regs_13_6 <= _T_2405;
    end
    if (io_load) begin
      regs_13_7 <= io_data[215];
    end else if (_T_2413) begin
      regs_13_7 <= 1'h0;
    end else if (!(_T_2414)) begin
      regs_13_7 <= _T_2415;
    end
    if (io_load) begin
      regs_13_8 <= io_data[216];
    end else if (_T_2423) begin
      regs_13_8 <= 1'h0;
    end else if (!(_T_2424)) begin
      regs_13_8 <= _T_2425;
    end
    if (io_load) begin
      regs_13_9 <= io_data[217];
    end else if (_T_2433) begin
      regs_13_9 <= 1'h0;
    end else if (!(_T_2434)) begin
      regs_13_9 <= _T_2435;
    end
    if (io_load) begin
      regs_13_10 <= io_data[218];
    end else if (_T_2443) begin
      regs_13_10 <= 1'h0;
    end else if (!(_T_2444)) begin
      regs_13_10 <= _T_2445;
    end
    if (io_load) begin
      regs_13_11 <= io_data[219];
    end else if (_T_2453) begin
      regs_13_11 <= 1'h0;
    end else if (!(_T_2454)) begin
      regs_13_11 <= _T_2455;
    end
    if (io_load) begin
      regs_13_12 <= io_data[220];
    end else if (_T_2463) begin
      regs_13_12 <= 1'h0;
    end else if (!(_T_2464)) begin
      regs_13_12 <= _T_2465;
    end
    if (io_load) begin
      regs_13_13 <= io_data[221];
    end else if (_T_2473) begin
      regs_13_13 <= 1'h0;
    end else if (!(_T_2474)) begin
      regs_13_13 <= _T_2475;
    end
    if (io_load) begin
      regs_13_14 <= io_data[222];
    end else if (_T_2483) begin
      regs_13_14 <= 1'h0;
    end else if (!(_T_2484)) begin
      regs_13_14 <= _T_2485;
    end
    if (io_load) begin
      regs_13_15 <= io_data[223];
    end else if (_T_2493) begin
      regs_13_15 <= 1'h0;
    end else if (!(_T_2494)) begin
      regs_13_15 <= _T_2495;
    end
    if (io_load) begin
      regs_14_0 <= io_data[224];
    end else if (_T_2503) begin
      regs_14_0 <= 1'h0;
    end else if (!(_T_2504)) begin
      regs_14_0 <= _T_2505;
    end
    if (io_load) begin
      regs_14_1 <= io_data[225];
    end else if (_T_2513) begin
      regs_14_1 <= 1'h0;
    end else if (!(_T_2514)) begin
      regs_14_1 <= _T_2515;
    end
    if (io_load) begin
      regs_14_2 <= io_data[226];
    end else if (_T_2523) begin
      regs_14_2 <= 1'h0;
    end else if (!(_T_2524)) begin
      regs_14_2 <= _T_2525;
    end
    if (io_load) begin
      regs_14_3 <= io_data[227];
    end else if (_T_2533) begin
      regs_14_3 <= 1'h0;
    end else if (!(_T_2534)) begin
      regs_14_3 <= _T_2535;
    end
    if (io_load) begin
      regs_14_4 <= io_data[228];
    end else if (_T_2543) begin
      regs_14_4 <= 1'h0;
    end else if (!(_T_2544)) begin
      regs_14_4 <= _T_2545;
    end
    if (io_load) begin
      regs_14_5 <= io_data[229];
    end else if (_T_2553) begin
      regs_14_5 <= 1'h0;
    end else if (!(_T_2554)) begin
      regs_14_5 <= _T_2555;
    end
    if (io_load) begin
      regs_14_6 <= io_data[230];
    end else if (_T_2563) begin
      regs_14_6 <= 1'h0;
    end else if (!(_T_2564)) begin
      regs_14_6 <= _T_2565;
    end
    if (io_load) begin
      regs_14_7 <= io_data[231];
    end else if (_T_2573) begin
      regs_14_7 <= 1'h0;
    end else if (!(_T_2574)) begin
      regs_14_7 <= _T_2575;
    end
    if (io_load) begin
      regs_14_8 <= io_data[232];
    end else if (_T_2583) begin
      regs_14_8 <= 1'h0;
    end else if (!(_T_2584)) begin
      regs_14_8 <= _T_2585;
    end
    if (io_load) begin
      regs_14_9 <= io_data[233];
    end else if (_T_2593) begin
      regs_14_9 <= 1'h0;
    end else if (!(_T_2594)) begin
      regs_14_9 <= _T_2595;
    end
    if (io_load) begin
      regs_14_10 <= io_data[234];
    end else if (_T_2603) begin
      regs_14_10 <= 1'h0;
    end else if (!(_T_2604)) begin
      regs_14_10 <= _T_2605;
    end
    if (io_load) begin
      regs_14_11 <= io_data[235];
    end else if (_T_2613) begin
      regs_14_11 <= 1'h0;
    end else if (!(_T_2614)) begin
      regs_14_11 <= _T_2615;
    end
    if (io_load) begin
      regs_14_12 <= io_data[236];
    end else if (_T_2623) begin
      regs_14_12 <= 1'h0;
    end else if (!(_T_2624)) begin
      regs_14_12 <= _T_2625;
    end
    if (io_load) begin
      regs_14_13 <= io_data[237];
    end else if (_T_2633) begin
      regs_14_13 <= 1'h0;
    end else if (!(_T_2634)) begin
      regs_14_13 <= _T_2635;
    end
    if (io_load) begin
      regs_14_14 <= io_data[238];
    end else if (_T_2643) begin
      regs_14_14 <= 1'h0;
    end else if (!(_T_2644)) begin
      regs_14_14 <= _T_2645;
    end
    if (io_load) begin
      regs_14_15 <= io_data[239];
    end else if (_T_2653) begin
      regs_14_15 <= 1'h0;
    end else if (!(_T_2654)) begin
      regs_14_15 <= _T_2655;
    end
    if (io_load) begin
      regs_15_0 <= io_data[240];
    end else if (_T_2663) begin
      regs_15_0 <= 1'h0;
    end else if (!(_T_2664)) begin
      regs_15_0 <= _T_2665;
    end
    if (io_load) begin
      regs_15_1 <= io_data[241];
    end else if (_T_2673) begin
      regs_15_1 <= 1'h0;
    end else if (!(_T_2674)) begin
      regs_15_1 <= _T_2675;
    end
    if (io_load) begin
      regs_15_2 <= io_data[242];
    end else if (_T_2683) begin
      regs_15_2 <= 1'h0;
    end else if (!(_T_2684)) begin
      regs_15_2 <= _T_2685;
    end
    if (io_load) begin
      regs_15_3 <= io_data[243];
    end else if (_T_2693) begin
      regs_15_3 <= 1'h0;
    end else if (!(_T_2694)) begin
      regs_15_3 <= _T_2695;
    end
    if (io_load) begin
      regs_15_4 <= io_data[244];
    end else if (_T_2703) begin
      regs_15_4 <= 1'h0;
    end else if (!(_T_2704)) begin
      regs_15_4 <= _T_2705;
    end
    if (io_load) begin
      regs_15_5 <= io_data[245];
    end else if (_T_2713) begin
      regs_15_5 <= 1'h0;
    end else if (!(_T_2714)) begin
      regs_15_5 <= _T_2715;
    end
    if (io_load) begin
      regs_15_6 <= io_data[246];
    end else if (_T_2723) begin
      regs_15_6 <= 1'h0;
    end else if (!(_T_2724)) begin
      regs_15_6 <= _T_2725;
    end
    if (io_load) begin
      regs_15_7 <= io_data[247];
    end else if (_T_2733) begin
      regs_15_7 <= 1'h0;
    end else if (!(_T_2734)) begin
      regs_15_7 <= _T_2735;
    end
    if (io_load) begin
      regs_15_8 <= io_data[248];
    end else if (_T_2743) begin
      regs_15_8 <= 1'h0;
    end else if (!(_T_2744)) begin
      regs_15_8 <= _T_2745;
    end
    if (io_load) begin
      regs_15_9 <= io_data[249];
    end else if (_T_2753) begin
      regs_15_9 <= 1'h0;
    end else if (!(_T_2754)) begin
      regs_15_9 <= _T_2755;
    end
    if (io_load) begin
      regs_15_10 <= io_data[250];
    end else if (_T_2763) begin
      regs_15_10 <= 1'h0;
    end else if (!(_T_2764)) begin
      regs_15_10 <= _T_2765;
    end
    if (io_load) begin
      regs_15_11 <= io_data[251];
    end else if (_T_2773) begin
      regs_15_11 <= 1'h0;
    end else if (!(_T_2774)) begin
      regs_15_11 <= _T_2775;
    end
    if (io_load) begin
      regs_15_12 <= io_data[252];
    end else if (_T_2783) begin
      regs_15_12 <= 1'h0;
    end else if (!(_T_2784)) begin
      regs_15_12 <= _T_2785;
    end
    if (io_load) begin
      regs_15_13 <= io_data[253];
    end else if (_T_2793) begin
      regs_15_13 <= 1'h0;
    end else if (!(_T_2794)) begin
      regs_15_13 <= _T_2795;
    end
    if (io_load) begin
      regs_15_14 <= io_data[254];
    end else if (_T_2803) begin
      regs_15_14 <= 1'h0;
    end else if (!(_T_2804)) begin
      regs_15_14 <= _T_2805;
    end
    if (io_load) begin
      regs_15_15 <= io_data[255];
    end else if (_T_2813) begin
      regs_15_15 <= 1'h0;
    end else if (!(_T_2814)) begin
      regs_15_15 <= _T_2815;
    end
  end
endmodule
