module ConwaylifeBetter(
  input          clock,
  input          reset,
  input          io_load,
  input  [255:0] io_data,
  output [255:0] io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] regs; // @[ConwaylifeBetter.scala 10:17]
  wire [1:0] _T_265 = regs[255] + regs[240]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_513 = {{1'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_266 = _T_265 + _GEN_513; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_514 = {{2'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_267 = _T_266 + _GEN_514; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_515 = {{3'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_268 = _T_267 + _GEN_515; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_516 = {{4'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_269 = _T_268 + _GEN_516; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_517 = {{5'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_270 = _T_269 + _GEN_517; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_518 = {{6'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_271 = _T_270 + _GEN_518; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_272 = 8'h2 == _T_271; // @[Conditional.scala 37:30]
  wire  _T_274 = 8'h3 == _T_271; // @[Conditional.scala 37:30]
  wire  _GEN_1 = _T_272 ? regs[0] : _T_274; // @[Conditional.scala 40:58]
  wire [1:0] _T_283 = regs[240] + regs[241]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_519 = {{1'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_284 = _T_283 + _GEN_519; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_520 = {{2'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_285 = _T_284 + _GEN_520; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_521 = {{3'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_286 = _T_285 + _GEN_521; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_522 = {{4'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_287 = _T_286 + _GEN_522; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_523 = {{5'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_288 = _T_287 + _GEN_523; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_524 = {{6'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_289 = _T_288 + _GEN_524; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_290 = 8'h2 == _T_289; // @[Conditional.scala 37:30]
  wire  _T_292 = 8'h3 == _T_289; // @[Conditional.scala 37:30]
  wire  _GEN_3 = _T_290 ? regs[1] : _T_292; // @[Conditional.scala 40:58]
  wire [1:0] _T_301 = regs[241] + regs[242]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_525 = {{1'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_302 = _T_301 + _GEN_525; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_526 = {{2'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_303 = _T_302 + _GEN_526; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_527 = {{3'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_304 = _T_303 + _GEN_527; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_528 = {{4'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_305 = _T_304 + _GEN_528; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_529 = {{5'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_306 = _T_305 + _GEN_529; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_530 = {{6'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_307 = _T_306 + _GEN_530; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_308 = 8'h2 == _T_307; // @[Conditional.scala 37:30]
  wire  _T_310 = 8'h3 == _T_307; // @[Conditional.scala 37:30]
  wire  _GEN_5 = _T_308 ? regs[2] : _T_310; // @[Conditional.scala 40:58]
  wire [1:0] _T_319 = regs[242] + regs[243]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_531 = {{1'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_320 = _T_319 + _GEN_531; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_532 = {{2'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_321 = _T_320 + _GEN_532; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_533 = {{3'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_322 = _T_321 + _GEN_533; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_534 = {{4'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_323 = _T_322 + _GEN_534; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_535 = {{5'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_324 = _T_323 + _GEN_535; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_536 = {{6'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_325 = _T_324 + _GEN_536; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_326 = 8'h2 == _T_325; // @[Conditional.scala 37:30]
  wire  _T_328 = 8'h3 == _T_325; // @[Conditional.scala 37:30]
  wire  _GEN_7 = _T_326 ? regs[3] : _T_328; // @[Conditional.scala 40:58]
  wire [1:0] _T_337 = regs[243] + regs[244]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_537 = {{1'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_338 = _T_337 + _GEN_537; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_538 = {{2'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_339 = _T_338 + _GEN_538; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_539 = {{3'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_340 = _T_339 + _GEN_539; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_540 = {{4'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_341 = _T_340 + _GEN_540; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_541 = {{5'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_342 = _T_341 + _GEN_541; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_542 = {{6'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_343 = _T_342 + _GEN_542; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_344 = 8'h2 == _T_343; // @[Conditional.scala 37:30]
  wire  _T_346 = 8'h3 == _T_343; // @[Conditional.scala 37:30]
  wire  _GEN_9 = _T_344 ? regs[4] : _T_346; // @[Conditional.scala 40:58]
  wire [1:0] _T_355 = regs[244] + regs[245]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_543 = {{1'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_356 = _T_355 + _GEN_543; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_544 = {{2'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_357 = _T_356 + _GEN_544; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_545 = {{3'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_358 = _T_357 + _GEN_545; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_546 = {{4'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_359 = _T_358 + _GEN_546; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_547 = {{5'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_360 = _T_359 + _GEN_547; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_548 = {{6'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_361 = _T_360 + _GEN_548; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_362 = 8'h2 == _T_361; // @[Conditional.scala 37:30]
  wire  _T_364 = 8'h3 == _T_361; // @[Conditional.scala 37:30]
  wire  _GEN_11 = _T_362 ? regs[5] : _T_364; // @[Conditional.scala 40:58]
  wire [1:0] _T_373 = regs[245] + regs[246]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_549 = {{1'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_374 = _T_373 + _GEN_549; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_550 = {{2'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_375 = _T_374 + _GEN_550; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_551 = {{3'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_376 = _T_375 + _GEN_551; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_552 = {{4'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_377 = _T_376 + _GEN_552; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_553 = {{5'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_378 = _T_377 + _GEN_553; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_554 = {{6'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_379 = _T_378 + _GEN_554; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_380 = 8'h2 == _T_379; // @[Conditional.scala 37:30]
  wire  _T_382 = 8'h3 == _T_379; // @[Conditional.scala 37:30]
  wire  _GEN_13 = _T_380 ? regs[6] : _T_382; // @[Conditional.scala 40:58]
  wire [1:0] _T_391 = regs[246] + regs[247]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_555 = {{1'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_392 = _T_391 + _GEN_555; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_556 = {{2'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_393 = _T_392 + _GEN_556; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_557 = {{3'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_394 = _T_393 + _GEN_557; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_558 = {{4'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_395 = _T_394 + _GEN_558; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_559 = {{5'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_396 = _T_395 + _GEN_559; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_560 = {{6'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_397 = _T_396 + _GEN_560; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_398 = 8'h2 == _T_397; // @[Conditional.scala 37:30]
  wire  _T_400 = 8'h3 == _T_397; // @[Conditional.scala 37:30]
  wire  _GEN_15 = _T_398 ? regs[7] : _T_400; // @[Conditional.scala 40:58]
  wire [1:0] _T_409 = regs[247] + regs[248]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_561 = {{1'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_410 = _T_409 + _GEN_561; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_562 = {{2'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_411 = _T_410 + _GEN_562; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_563 = {{3'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_412 = _T_411 + _GEN_563; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_564 = {{4'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_413 = _T_412 + _GEN_564; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_565 = {{5'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_414 = _T_413 + _GEN_565; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_566 = {{6'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_415 = _T_414 + _GEN_566; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_416 = 8'h2 == _T_415; // @[Conditional.scala 37:30]
  wire  _T_418 = 8'h3 == _T_415; // @[Conditional.scala 37:30]
  wire  _GEN_17 = _T_416 ? regs[8] : _T_418; // @[Conditional.scala 40:58]
  wire [1:0] _T_427 = regs[248] + regs[249]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_567 = {{1'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_428 = _T_427 + _GEN_567; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_568 = {{2'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_429 = _T_428 + _GEN_568; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_569 = {{3'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_430 = _T_429 + _GEN_569; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_570 = {{4'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_431 = _T_430 + _GEN_570; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_571 = {{5'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_432 = _T_431 + _GEN_571; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_572 = {{6'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_433 = _T_432 + _GEN_572; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_434 = 8'h2 == _T_433; // @[Conditional.scala 37:30]
  wire  _T_436 = 8'h3 == _T_433; // @[Conditional.scala 37:30]
  wire  _GEN_19 = _T_434 ? regs[9] : _T_436; // @[Conditional.scala 40:58]
  wire [1:0] _T_445 = regs[249] + regs[250]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_573 = {{1'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_446 = _T_445 + _GEN_573; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_574 = {{2'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_447 = _T_446 + _GEN_574; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_575 = {{3'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_448 = _T_447 + _GEN_575; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_576 = {{4'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_449 = _T_448 + _GEN_576; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_577 = {{5'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_450 = _T_449 + _GEN_577; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_578 = {{6'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_451 = _T_450 + _GEN_578; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_452 = 8'h2 == _T_451; // @[Conditional.scala 37:30]
  wire  _T_454 = 8'h3 == _T_451; // @[Conditional.scala 37:30]
  wire  _GEN_21 = _T_452 ? regs[10] : _T_454; // @[Conditional.scala 40:58]
  wire [1:0] _T_463 = regs[250] + regs[251]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_579 = {{1'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_464 = _T_463 + _GEN_579; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_580 = {{2'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_465 = _T_464 + _GEN_580; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_581 = {{3'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_466 = _T_465 + _GEN_581; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_582 = {{4'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_467 = _T_466 + _GEN_582; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_583 = {{5'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_468 = _T_467 + _GEN_583; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_584 = {{6'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_469 = _T_468 + _GEN_584; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_470 = 8'h2 == _T_469; // @[Conditional.scala 37:30]
  wire  _T_472 = 8'h3 == _T_469; // @[Conditional.scala 37:30]
  wire  _GEN_23 = _T_470 ? regs[11] : _T_472; // @[Conditional.scala 40:58]
  wire [1:0] _T_481 = regs[251] + regs[252]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_585 = {{1'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_482 = _T_481 + _GEN_585; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_586 = {{2'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_483 = _T_482 + _GEN_586; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_587 = {{3'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_484 = _T_483 + _GEN_587; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_588 = {{4'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_485 = _T_484 + _GEN_588; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_589 = {{5'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_486 = _T_485 + _GEN_589; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_590 = {{6'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_487 = _T_486 + _GEN_590; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_488 = 8'h2 == _T_487; // @[Conditional.scala 37:30]
  wire  _T_490 = 8'h3 == _T_487; // @[Conditional.scala 37:30]
  wire  _GEN_25 = _T_488 ? regs[12] : _T_490; // @[Conditional.scala 40:58]
  wire [1:0] _T_499 = regs[252] + regs[253]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_591 = {{1'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_500 = _T_499 + _GEN_591; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_592 = {{2'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_501 = _T_500 + _GEN_592; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_593 = {{3'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_502 = _T_501 + _GEN_593; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_594 = {{4'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_503 = _T_502 + _GEN_594; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_595 = {{5'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_504 = _T_503 + _GEN_595; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_596 = {{6'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_505 = _T_504 + _GEN_596; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_506 = 8'h2 == _T_505; // @[Conditional.scala 37:30]
  wire  _T_508 = 8'h3 == _T_505; // @[Conditional.scala 37:30]
  wire  _GEN_27 = _T_506 ? regs[13] : _T_508; // @[Conditional.scala 40:58]
  wire [1:0] _T_517 = regs[253] + regs[254]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_597 = {{1'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_518 = _T_517 + _GEN_597; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_598 = {{2'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_519 = _T_518 + _GEN_598; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_599 = {{3'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_520 = _T_519 + _GEN_599; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_600 = {{4'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_521 = _T_520 + _GEN_600; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_601 = {{5'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_522 = _T_521 + _GEN_601; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_602 = {{6'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_523 = _T_522 + _GEN_602; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_524 = 8'h2 == _T_523; // @[Conditional.scala 37:30]
  wire  _T_526 = 8'h3 == _T_523; // @[Conditional.scala 37:30]
  wire  _GEN_29 = _T_524 ? regs[14] : _T_526; // @[Conditional.scala 40:58]
  wire [1:0] _T_535 = regs[254] + regs[255]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_603 = {{1'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_536 = _T_535 + _GEN_603; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_604 = {{2'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_537 = _T_536 + _GEN_604; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_605 = {{3'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_538 = _T_537 + _GEN_605; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_606 = {{4'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_539 = _T_538 + _GEN_606; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_607 = {{5'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_540 = _T_539 + _GEN_607; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_608 = {{6'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_541 = _T_540 + _GEN_608; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_542 = 8'h2 == _T_541; // @[Conditional.scala 37:30]
  wire  _T_544 = 8'h3 == _T_541; // @[Conditional.scala 37:30]
  wire  _GEN_31 = _T_542 ? regs[15] : _T_544; // @[Conditional.scala 40:58]
  wire [1:0] _T_553 = regs[15] + regs[0]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_609 = {{1'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_554 = _T_553 + _GEN_609; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_610 = {{2'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_555 = _T_554 + _GEN_610; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_611 = {{3'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_556 = _T_555 + _GEN_611; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_612 = {{4'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_557 = _T_556 + _GEN_612; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_613 = {{5'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_558 = _T_557 + _GEN_613; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_614 = {{6'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_559 = _T_558 + _GEN_614; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_560 = 8'h2 == _T_559; // @[Conditional.scala 37:30]
  wire  _T_562 = 8'h3 == _T_559; // @[Conditional.scala 37:30]
  wire  _GEN_33 = _T_560 ? regs[16] : _T_562; // @[Conditional.scala 40:58]
  wire [1:0] _T_571 = regs[0] + regs[1]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_615 = {{1'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_572 = _T_571 + _GEN_615; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_616 = {{2'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_573 = _T_572 + _GEN_616; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_617 = {{3'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_574 = _T_573 + _GEN_617; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_618 = {{4'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_575 = _T_574 + _GEN_618; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_619 = {{5'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_576 = _T_575 + _GEN_619; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_620 = {{6'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_577 = _T_576 + _GEN_620; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_578 = 8'h2 == _T_577; // @[Conditional.scala 37:30]
  wire  _T_580 = 8'h3 == _T_577; // @[Conditional.scala 37:30]
  wire  _GEN_35 = _T_578 ? regs[17] : _T_580; // @[Conditional.scala 40:58]
  wire [1:0] _T_589 = regs[1] + regs[2]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_621 = {{1'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_590 = _T_589 + _GEN_621; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_622 = {{2'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_591 = _T_590 + _GEN_622; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_623 = {{3'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_592 = _T_591 + _GEN_623; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_624 = {{4'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_593 = _T_592 + _GEN_624; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_625 = {{5'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_594 = _T_593 + _GEN_625; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_626 = {{6'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_595 = _T_594 + _GEN_626; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_596 = 8'h2 == _T_595; // @[Conditional.scala 37:30]
  wire  _T_598 = 8'h3 == _T_595; // @[Conditional.scala 37:30]
  wire  _GEN_37 = _T_596 ? regs[18] : _T_598; // @[Conditional.scala 40:58]
  wire [1:0] _T_607 = regs[2] + regs[3]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_627 = {{1'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_608 = _T_607 + _GEN_627; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_628 = {{2'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_609 = _T_608 + _GEN_628; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_629 = {{3'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_610 = _T_609 + _GEN_629; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_630 = {{4'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_611 = _T_610 + _GEN_630; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_631 = {{5'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_612 = _T_611 + _GEN_631; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_632 = {{6'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_613 = _T_612 + _GEN_632; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_614 = 8'h2 == _T_613; // @[Conditional.scala 37:30]
  wire  _T_616 = 8'h3 == _T_613; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_614 ? regs[19] : _T_616; // @[Conditional.scala 40:58]
  wire [1:0] _T_625 = regs[3] + regs[4]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_633 = {{1'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_626 = _T_625 + _GEN_633; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_634 = {{2'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_627 = _T_626 + _GEN_634; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_635 = {{3'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_628 = _T_627 + _GEN_635; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_636 = {{4'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_629 = _T_628 + _GEN_636; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_637 = {{5'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_630 = _T_629 + _GEN_637; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_638 = {{6'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_631 = _T_630 + _GEN_638; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_632 = 8'h2 == _T_631; // @[Conditional.scala 37:30]
  wire  _T_634 = 8'h3 == _T_631; // @[Conditional.scala 37:30]
  wire  _GEN_41 = _T_632 ? regs[20] : _T_634; // @[Conditional.scala 40:58]
  wire [1:0] _T_643 = regs[4] + regs[5]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_639 = {{1'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_644 = _T_643 + _GEN_639; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_640 = {{2'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_645 = _T_644 + _GEN_640; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_641 = {{3'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_646 = _T_645 + _GEN_641; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_642 = {{4'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_647 = _T_646 + _GEN_642; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_643 = {{5'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_648 = _T_647 + _GEN_643; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_644 = {{6'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_649 = _T_648 + _GEN_644; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_650 = 8'h2 == _T_649; // @[Conditional.scala 37:30]
  wire  _T_652 = 8'h3 == _T_649; // @[Conditional.scala 37:30]
  wire  _GEN_43 = _T_650 ? regs[21] : _T_652; // @[Conditional.scala 40:58]
  wire [1:0] _T_661 = regs[5] + regs[6]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_645 = {{1'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_662 = _T_661 + _GEN_645; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_646 = {{2'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_663 = _T_662 + _GEN_646; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_647 = {{3'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_664 = _T_663 + _GEN_647; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_648 = {{4'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_665 = _T_664 + _GEN_648; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_649 = {{5'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_666 = _T_665 + _GEN_649; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_650 = {{6'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_667 = _T_666 + _GEN_650; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_668 = 8'h2 == _T_667; // @[Conditional.scala 37:30]
  wire  _T_670 = 8'h3 == _T_667; // @[Conditional.scala 37:30]
  wire  _GEN_45 = _T_668 ? regs[22] : _T_670; // @[Conditional.scala 40:58]
  wire [1:0] _T_679 = regs[6] + regs[7]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_651 = {{1'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_680 = _T_679 + _GEN_651; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_652 = {{2'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_681 = _T_680 + _GEN_652; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_653 = {{3'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_682 = _T_681 + _GEN_653; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_654 = {{4'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_683 = _T_682 + _GEN_654; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_655 = {{5'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_684 = _T_683 + _GEN_655; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_656 = {{6'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_685 = _T_684 + _GEN_656; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_686 = 8'h2 == _T_685; // @[Conditional.scala 37:30]
  wire  _T_688 = 8'h3 == _T_685; // @[Conditional.scala 37:30]
  wire  _GEN_47 = _T_686 ? regs[23] : _T_688; // @[Conditional.scala 40:58]
  wire [1:0] _T_697 = regs[7] + regs[8]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_657 = {{1'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_698 = _T_697 + _GEN_657; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_658 = {{2'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_699 = _T_698 + _GEN_658; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_659 = {{3'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_700 = _T_699 + _GEN_659; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_660 = {{4'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_701 = _T_700 + _GEN_660; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_661 = {{5'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_702 = _T_701 + _GEN_661; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_662 = {{6'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_703 = _T_702 + _GEN_662; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_704 = 8'h2 == _T_703; // @[Conditional.scala 37:30]
  wire  _T_706 = 8'h3 == _T_703; // @[Conditional.scala 37:30]
  wire  _GEN_49 = _T_704 ? regs[24] : _T_706; // @[Conditional.scala 40:58]
  wire [1:0] _T_715 = regs[8] + regs[9]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_663 = {{1'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_716 = _T_715 + _GEN_663; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_664 = {{2'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_717 = _T_716 + _GEN_664; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_665 = {{3'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_718 = _T_717 + _GEN_665; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_666 = {{4'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_719 = _T_718 + _GEN_666; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_667 = {{5'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_720 = _T_719 + _GEN_667; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_668 = {{6'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_721 = _T_720 + _GEN_668; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_722 = 8'h2 == _T_721; // @[Conditional.scala 37:30]
  wire  _T_724 = 8'h3 == _T_721; // @[Conditional.scala 37:30]
  wire  _GEN_51 = _T_722 ? regs[25] : _T_724; // @[Conditional.scala 40:58]
  wire [1:0] _T_733 = regs[9] + regs[10]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_669 = {{1'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_734 = _T_733 + _GEN_669; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_670 = {{2'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_735 = _T_734 + _GEN_670; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_671 = {{3'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_736 = _T_735 + _GEN_671; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_672 = {{4'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_737 = _T_736 + _GEN_672; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_673 = {{5'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_738 = _T_737 + _GEN_673; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_674 = {{6'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_739 = _T_738 + _GEN_674; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_740 = 8'h2 == _T_739; // @[Conditional.scala 37:30]
  wire  _T_742 = 8'h3 == _T_739; // @[Conditional.scala 37:30]
  wire  _GEN_53 = _T_740 ? regs[26] : _T_742; // @[Conditional.scala 40:58]
  wire [1:0] _T_751 = regs[10] + regs[11]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_675 = {{1'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_752 = _T_751 + _GEN_675; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_676 = {{2'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_753 = _T_752 + _GEN_676; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_677 = {{3'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_754 = _T_753 + _GEN_677; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_678 = {{4'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_755 = _T_754 + _GEN_678; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_679 = {{5'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_756 = _T_755 + _GEN_679; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_680 = {{6'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_757 = _T_756 + _GEN_680; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_758 = 8'h2 == _T_757; // @[Conditional.scala 37:30]
  wire  _T_760 = 8'h3 == _T_757; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_758 ? regs[27] : _T_760; // @[Conditional.scala 40:58]
  wire [1:0] _T_769 = regs[11] + regs[12]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_681 = {{1'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_770 = _T_769 + _GEN_681; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_682 = {{2'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_771 = _T_770 + _GEN_682; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_683 = {{3'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_772 = _T_771 + _GEN_683; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_684 = {{4'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_773 = _T_772 + _GEN_684; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_685 = {{5'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_774 = _T_773 + _GEN_685; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_686 = {{6'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_775 = _T_774 + _GEN_686; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_776 = 8'h2 == _T_775; // @[Conditional.scala 37:30]
  wire  _T_778 = 8'h3 == _T_775; // @[Conditional.scala 37:30]
  wire  _GEN_57 = _T_776 ? regs[28] : _T_778; // @[Conditional.scala 40:58]
  wire [1:0] _T_787 = regs[12] + regs[13]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_687 = {{1'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_788 = _T_787 + _GEN_687; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_688 = {{2'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_789 = _T_788 + _GEN_688; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_689 = {{3'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_790 = _T_789 + _GEN_689; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_690 = {{4'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_791 = _T_790 + _GEN_690; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_691 = {{5'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_792 = _T_791 + _GEN_691; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_692 = {{6'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_793 = _T_792 + _GEN_692; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_794 = 8'h2 == _T_793; // @[Conditional.scala 37:30]
  wire  _T_796 = 8'h3 == _T_793; // @[Conditional.scala 37:30]
  wire  _GEN_59 = _T_794 ? regs[29] : _T_796; // @[Conditional.scala 40:58]
  wire [1:0] _T_805 = regs[13] + regs[14]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_693 = {{1'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_806 = _T_805 + _GEN_693; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_694 = {{2'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_807 = _T_806 + _GEN_694; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_695 = {{3'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_808 = _T_807 + _GEN_695; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_696 = {{4'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_809 = _T_808 + _GEN_696; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_697 = {{5'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_810 = _T_809 + _GEN_697; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_698 = {{6'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_811 = _T_810 + _GEN_698; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_812 = 8'h2 == _T_811; // @[Conditional.scala 37:30]
  wire  _T_814 = 8'h3 == _T_811; // @[Conditional.scala 37:30]
  wire  _GEN_61 = _T_812 ? regs[30] : _T_814; // @[Conditional.scala 40:58]
  wire [1:0] _T_823 = regs[14] + regs[15]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_699 = {{1'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_824 = _T_823 + _GEN_699; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_700 = {{2'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_825 = _T_824 + _GEN_700; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_701 = {{3'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_826 = _T_825 + _GEN_701; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_702 = {{4'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_827 = _T_826 + _GEN_702; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_703 = {{5'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_828 = _T_827 + _GEN_703; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_704 = {{6'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_829 = _T_828 + _GEN_704; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_830 = 8'h2 == _T_829; // @[Conditional.scala 37:30]
  wire  _T_832 = 8'h3 == _T_829; // @[Conditional.scala 37:30]
  wire  _GEN_63 = _T_830 ? regs[31] : _T_832; // @[Conditional.scala 40:58]
  wire [1:0] _T_841 = regs[31] + regs[16]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_705 = {{1'd0}, regs[17]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_842 = _T_841 + _GEN_705; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_706 = {{2'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_843 = _T_842 + _GEN_706; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_707 = {{3'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_844 = _T_843 + _GEN_707; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_708 = {{4'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_845 = _T_844 + _GEN_708; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_709 = {{5'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_846 = _T_845 + _GEN_709; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_710 = {{6'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_847 = _T_846 + _GEN_710; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_848 = 8'h2 == _T_847; // @[Conditional.scala 37:30]
  wire  _T_850 = 8'h3 == _T_847; // @[Conditional.scala 37:30]
  wire  _GEN_65 = _T_848 ? regs[32] : _T_850; // @[Conditional.scala 40:58]
  wire [1:0] _T_859 = regs[16] + regs[17]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_711 = {{1'd0}, regs[18]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_860 = _T_859 + _GEN_711; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_712 = {{2'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_861 = _T_860 + _GEN_712; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_713 = {{3'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_862 = _T_861 + _GEN_713; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_714 = {{4'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_863 = _T_862 + _GEN_714; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_715 = {{5'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_864 = _T_863 + _GEN_715; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_716 = {{6'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_865 = _T_864 + _GEN_716; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_866 = 8'h2 == _T_865; // @[Conditional.scala 37:30]
  wire  _T_868 = 8'h3 == _T_865; // @[Conditional.scala 37:30]
  wire  _GEN_67 = _T_866 ? regs[33] : _T_868; // @[Conditional.scala 40:58]
  wire [1:0] _T_877 = regs[17] + regs[18]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_717 = {{1'd0}, regs[19]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_878 = _T_877 + _GEN_717; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_718 = {{2'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_879 = _T_878 + _GEN_718; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_719 = {{3'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_880 = _T_879 + _GEN_719; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_720 = {{4'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_881 = _T_880 + _GEN_720; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_721 = {{5'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_882 = _T_881 + _GEN_721; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_722 = {{6'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_883 = _T_882 + _GEN_722; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_884 = 8'h2 == _T_883; // @[Conditional.scala 37:30]
  wire  _T_886 = 8'h3 == _T_883; // @[Conditional.scala 37:30]
  wire  _GEN_69 = _T_884 ? regs[34] : _T_886; // @[Conditional.scala 40:58]
  wire [1:0] _T_895 = regs[18] + regs[19]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_723 = {{1'd0}, regs[20]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_896 = _T_895 + _GEN_723; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_724 = {{2'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_897 = _T_896 + _GEN_724; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_725 = {{3'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_898 = _T_897 + _GEN_725; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_726 = {{4'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_899 = _T_898 + _GEN_726; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_727 = {{5'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_900 = _T_899 + _GEN_727; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_728 = {{6'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_901 = _T_900 + _GEN_728; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_902 = 8'h2 == _T_901; // @[Conditional.scala 37:30]
  wire  _T_904 = 8'h3 == _T_901; // @[Conditional.scala 37:30]
  wire  _GEN_71 = _T_902 ? regs[35] : _T_904; // @[Conditional.scala 40:58]
  wire [1:0] _T_913 = regs[19] + regs[20]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_729 = {{1'd0}, regs[21]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_914 = _T_913 + _GEN_729; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_730 = {{2'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_915 = _T_914 + _GEN_730; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_731 = {{3'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_916 = _T_915 + _GEN_731; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_732 = {{4'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_917 = _T_916 + _GEN_732; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_733 = {{5'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_918 = _T_917 + _GEN_733; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_734 = {{6'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_919 = _T_918 + _GEN_734; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_920 = 8'h2 == _T_919; // @[Conditional.scala 37:30]
  wire  _T_922 = 8'h3 == _T_919; // @[Conditional.scala 37:30]
  wire  _GEN_73 = _T_920 ? regs[36] : _T_922; // @[Conditional.scala 40:58]
  wire [1:0] _T_931 = regs[20] + regs[21]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_735 = {{1'd0}, regs[22]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_932 = _T_931 + _GEN_735; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_736 = {{2'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_933 = _T_932 + _GEN_736; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_737 = {{3'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_934 = _T_933 + _GEN_737; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_738 = {{4'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_935 = _T_934 + _GEN_738; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_739 = {{5'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_936 = _T_935 + _GEN_739; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_740 = {{6'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_937 = _T_936 + _GEN_740; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_938 = 8'h2 == _T_937; // @[Conditional.scala 37:30]
  wire  _T_940 = 8'h3 == _T_937; // @[Conditional.scala 37:30]
  wire  _GEN_75 = _T_938 ? regs[37] : _T_940; // @[Conditional.scala 40:58]
  wire [1:0] _T_949 = regs[21] + regs[22]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_741 = {{1'd0}, regs[23]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_950 = _T_949 + _GEN_741; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_742 = {{2'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_951 = _T_950 + _GEN_742; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_743 = {{3'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_952 = _T_951 + _GEN_743; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_744 = {{4'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_953 = _T_952 + _GEN_744; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_745 = {{5'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_954 = _T_953 + _GEN_745; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_746 = {{6'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_955 = _T_954 + _GEN_746; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_956 = 8'h2 == _T_955; // @[Conditional.scala 37:30]
  wire  _T_958 = 8'h3 == _T_955; // @[Conditional.scala 37:30]
  wire  _GEN_77 = _T_956 ? regs[38] : _T_958; // @[Conditional.scala 40:58]
  wire [1:0] _T_967 = regs[22] + regs[23]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_747 = {{1'd0}, regs[24]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_968 = _T_967 + _GEN_747; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_748 = {{2'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_969 = _T_968 + _GEN_748; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_749 = {{3'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_970 = _T_969 + _GEN_749; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_750 = {{4'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_971 = _T_970 + _GEN_750; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_751 = {{5'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_972 = _T_971 + _GEN_751; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_752 = {{6'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_973 = _T_972 + _GEN_752; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_974 = 8'h2 == _T_973; // @[Conditional.scala 37:30]
  wire  _T_976 = 8'h3 == _T_973; // @[Conditional.scala 37:30]
  wire  _GEN_79 = _T_974 ? regs[39] : _T_976; // @[Conditional.scala 40:58]
  wire [1:0] _T_985 = regs[23] + regs[24]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_753 = {{1'd0}, regs[25]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_986 = _T_985 + _GEN_753; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_754 = {{2'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_987 = _T_986 + _GEN_754; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_755 = {{3'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_988 = _T_987 + _GEN_755; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_756 = {{4'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_989 = _T_988 + _GEN_756; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_757 = {{5'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_990 = _T_989 + _GEN_757; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_758 = {{6'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_991 = _T_990 + _GEN_758; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_992 = 8'h2 == _T_991; // @[Conditional.scala 37:30]
  wire  _T_994 = 8'h3 == _T_991; // @[Conditional.scala 37:30]
  wire  _GEN_81 = _T_992 ? regs[40] : _T_994; // @[Conditional.scala 40:58]
  wire [1:0] _T_1003 = regs[24] + regs[25]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_759 = {{1'd0}, regs[26]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1004 = _T_1003 + _GEN_759; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_760 = {{2'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1005 = _T_1004 + _GEN_760; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_761 = {{3'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1006 = _T_1005 + _GEN_761; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_762 = {{4'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1007 = _T_1006 + _GEN_762; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_763 = {{5'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1008 = _T_1007 + _GEN_763; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_764 = {{6'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1009 = _T_1008 + _GEN_764; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1010 = 8'h2 == _T_1009; // @[Conditional.scala 37:30]
  wire  _T_1012 = 8'h3 == _T_1009; // @[Conditional.scala 37:30]
  wire  _GEN_83 = _T_1010 ? regs[41] : _T_1012; // @[Conditional.scala 40:58]
  wire [1:0] _T_1021 = regs[25] + regs[26]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_765 = {{1'd0}, regs[27]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1022 = _T_1021 + _GEN_765; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_766 = {{2'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1023 = _T_1022 + _GEN_766; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_767 = {{3'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1024 = _T_1023 + _GEN_767; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_768 = {{4'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1025 = _T_1024 + _GEN_768; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_769 = {{5'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1026 = _T_1025 + _GEN_769; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_770 = {{6'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1027 = _T_1026 + _GEN_770; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1028 = 8'h2 == _T_1027; // @[Conditional.scala 37:30]
  wire  _T_1030 = 8'h3 == _T_1027; // @[Conditional.scala 37:30]
  wire  _GEN_85 = _T_1028 ? regs[42] : _T_1030; // @[Conditional.scala 40:58]
  wire [1:0] _T_1039 = regs[26] + regs[27]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_771 = {{1'd0}, regs[28]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1040 = _T_1039 + _GEN_771; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_772 = {{2'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1041 = _T_1040 + _GEN_772; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_773 = {{3'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1042 = _T_1041 + _GEN_773; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_774 = {{4'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1043 = _T_1042 + _GEN_774; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_775 = {{5'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1044 = _T_1043 + _GEN_775; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_776 = {{6'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1045 = _T_1044 + _GEN_776; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1046 = 8'h2 == _T_1045; // @[Conditional.scala 37:30]
  wire  _T_1048 = 8'h3 == _T_1045; // @[Conditional.scala 37:30]
  wire  _GEN_87 = _T_1046 ? regs[43] : _T_1048; // @[Conditional.scala 40:58]
  wire [1:0] _T_1057 = regs[27] + regs[28]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_777 = {{1'd0}, regs[29]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1058 = _T_1057 + _GEN_777; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_778 = {{2'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1059 = _T_1058 + _GEN_778; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_779 = {{3'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1060 = _T_1059 + _GEN_779; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_780 = {{4'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1061 = _T_1060 + _GEN_780; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_781 = {{5'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1062 = _T_1061 + _GEN_781; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_782 = {{6'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1063 = _T_1062 + _GEN_782; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1064 = 8'h2 == _T_1063; // @[Conditional.scala 37:30]
  wire  _T_1066 = 8'h3 == _T_1063; // @[Conditional.scala 37:30]
  wire  _GEN_89 = _T_1064 ? regs[44] : _T_1066; // @[Conditional.scala 40:58]
  wire [1:0] _T_1075 = regs[28] + regs[29]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_783 = {{1'd0}, regs[30]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1076 = _T_1075 + _GEN_783; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_784 = {{2'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1077 = _T_1076 + _GEN_784; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_785 = {{3'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1078 = _T_1077 + _GEN_785; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_786 = {{4'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1079 = _T_1078 + _GEN_786; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_787 = {{5'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1080 = _T_1079 + _GEN_787; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_788 = {{6'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1081 = _T_1080 + _GEN_788; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1082 = 8'h2 == _T_1081; // @[Conditional.scala 37:30]
  wire  _T_1084 = 8'h3 == _T_1081; // @[Conditional.scala 37:30]
  wire  _GEN_91 = _T_1082 ? regs[45] : _T_1084; // @[Conditional.scala 40:58]
  wire [1:0] _T_1093 = regs[29] + regs[30]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_789 = {{1'd0}, regs[31]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1094 = _T_1093 + _GEN_789; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_790 = {{2'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1095 = _T_1094 + _GEN_790; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_791 = {{3'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1096 = _T_1095 + _GEN_791; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_792 = {{4'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1097 = _T_1096 + _GEN_792; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_793 = {{5'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1098 = _T_1097 + _GEN_793; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_794 = {{6'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1099 = _T_1098 + _GEN_794; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1100 = 8'h2 == _T_1099; // @[Conditional.scala 37:30]
  wire  _T_1102 = 8'h3 == _T_1099; // @[Conditional.scala 37:30]
  wire  _GEN_93 = _T_1100 ? regs[46] : _T_1102; // @[Conditional.scala 40:58]
  wire [1:0] _T_1111 = regs[30] + regs[31]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_795 = {{1'd0}, regs[16]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1112 = _T_1111 + _GEN_795; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_796 = {{2'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1113 = _T_1112 + _GEN_796; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_797 = {{3'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1114 = _T_1113 + _GEN_797; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_798 = {{4'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1115 = _T_1114 + _GEN_798; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_799 = {{5'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1116 = _T_1115 + _GEN_799; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_800 = {{6'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1117 = _T_1116 + _GEN_800; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1118 = 8'h2 == _T_1117; // @[Conditional.scala 37:30]
  wire  _T_1120 = 8'h3 == _T_1117; // @[Conditional.scala 37:30]
  wire  _GEN_95 = _T_1118 ? regs[47] : _T_1120; // @[Conditional.scala 40:58]
  wire [1:0] _T_1129 = regs[47] + regs[32]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_801 = {{1'd0}, regs[33]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1130 = _T_1129 + _GEN_801; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_802 = {{2'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1131 = _T_1130 + _GEN_802; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_803 = {{3'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1132 = _T_1131 + _GEN_803; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_804 = {{4'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1133 = _T_1132 + _GEN_804; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_805 = {{5'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1134 = _T_1133 + _GEN_805; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_806 = {{6'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1135 = _T_1134 + _GEN_806; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1136 = 8'h2 == _T_1135; // @[Conditional.scala 37:30]
  wire  _T_1138 = 8'h3 == _T_1135; // @[Conditional.scala 37:30]
  wire  _GEN_97 = _T_1136 ? regs[48] : _T_1138; // @[Conditional.scala 40:58]
  wire [1:0] _T_1147 = regs[32] + regs[33]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_807 = {{1'd0}, regs[34]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1148 = _T_1147 + _GEN_807; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_808 = {{2'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1149 = _T_1148 + _GEN_808; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_809 = {{3'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1150 = _T_1149 + _GEN_809; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_810 = {{4'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1151 = _T_1150 + _GEN_810; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_811 = {{5'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1152 = _T_1151 + _GEN_811; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_812 = {{6'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1153 = _T_1152 + _GEN_812; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1154 = 8'h2 == _T_1153; // @[Conditional.scala 37:30]
  wire  _T_1156 = 8'h3 == _T_1153; // @[Conditional.scala 37:30]
  wire  _GEN_99 = _T_1154 ? regs[49] : _T_1156; // @[Conditional.scala 40:58]
  wire [1:0] _T_1165 = regs[33] + regs[34]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_813 = {{1'd0}, regs[35]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1166 = _T_1165 + _GEN_813; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_814 = {{2'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1167 = _T_1166 + _GEN_814; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_815 = {{3'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1168 = _T_1167 + _GEN_815; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_816 = {{4'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1169 = _T_1168 + _GEN_816; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_817 = {{5'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1170 = _T_1169 + _GEN_817; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_818 = {{6'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1171 = _T_1170 + _GEN_818; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1172 = 8'h2 == _T_1171; // @[Conditional.scala 37:30]
  wire  _T_1174 = 8'h3 == _T_1171; // @[Conditional.scala 37:30]
  wire  _GEN_101 = _T_1172 ? regs[50] : _T_1174; // @[Conditional.scala 40:58]
  wire [1:0] _T_1183 = regs[34] + regs[35]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_819 = {{1'd0}, regs[36]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1184 = _T_1183 + _GEN_819; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_820 = {{2'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1185 = _T_1184 + _GEN_820; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_821 = {{3'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1186 = _T_1185 + _GEN_821; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_822 = {{4'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1187 = _T_1186 + _GEN_822; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_823 = {{5'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1188 = _T_1187 + _GEN_823; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_824 = {{6'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1189 = _T_1188 + _GEN_824; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1190 = 8'h2 == _T_1189; // @[Conditional.scala 37:30]
  wire  _T_1192 = 8'h3 == _T_1189; // @[Conditional.scala 37:30]
  wire  _GEN_103 = _T_1190 ? regs[51] : _T_1192; // @[Conditional.scala 40:58]
  wire [1:0] _T_1201 = regs[35] + regs[36]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_825 = {{1'd0}, regs[37]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1202 = _T_1201 + _GEN_825; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_826 = {{2'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1203 = _T_1202 + _GEN_826; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_827 = {{3'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1204 = _T_1203 + _GEN_827; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_828 = {{4'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1205 = _T_1204 + _GEN_828; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_829 = {{5'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1206 = _T_1205 + _GEN_829; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_830 = {{6'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1207 = _T_1206 + _GEN_830; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1208 = 8'h2 == _T_1207; // @[Conditional.scala 37:30]
  wire  _T_1210 = 8'h3 == _T_1207; // @[Conditional.scala 37:30]
  wire  _GEN_105 = _T_1208 ? regs[52] : _T_1210; // @[Conditional.scala 40:58]
  wire [1:0] _T_1219 = regs[36] + regs[37]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_831 = {{1'd0}, regs[38]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1220 = _T_1219 + _GEN_831; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_832 = {{2'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1221 = _T_1220 + _GEN_832; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_833 = {{3'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1222 = _T_1221 + _GEN_833; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_834 = {{4'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1223 = _T_1222 + _GEN_834; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_835 = {{5'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1224 = _T_1223 + _GEN_835; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_836 = {{6'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1225 = _T_1224 + _GEN_836; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1226 = 8'h2 == _T_1225; // @[Conditional.scala 37:30]
  wire  _T_1228 = 8'h3 == _T_1225; // @[Conditional.scala 37:30]
  wire  _GEN_107 = _T_1226 ? regs[53] : _T_1228; // @[Conditional.scala 40:58]
  wire [1:0] _T_1237 = regs[37] + regs[38]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_837 = {{1'd0}, regs[39]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1238 = _T_1237 + _GEN_837; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_838 = {{2'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1239 = _T_1238 + _GEN_838; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_839 = {{3'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1240 = _T_1239 + _GEN_839; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_840 = {{4'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1241 = _T_1240 + _GEN_840; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_841 = {{5'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1242 = _T_1241 + _GEN_841; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_842 = {{6'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1243 = _T_1242 + _GEN_842; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1244 = 8'h2 == _T_1243; // @[Conditional.scala 37:30]
  wire  _T_1246 = 8'h3 == _T_1243; // @[Conditional.scala 37:30]
  wire  _GEN_109 = _T_1244 ? regs[54] : _T_1246; // @[Conditional.scala 40:58]
  wire [1:0] _T_1255 = regs[38] + regs[39]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_843 = {{1'd0}, regs[40]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1256 = _T_1255 + _GEN_843; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_844 = {{2'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1257 = _T_1256 + _GEN_844; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_845 = {{3'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1258 = _T_1257 + _GEN_845; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_846 = {{4'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1259 = _T_1258 + _GEN_846; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_847 = {{5'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1260 = _T_1259 + _GEN_847; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_848 = {{6'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1261 = _T_1260 + _GEN_848; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1262 = 8'h2 == _T_1261; // @[Conditional.scala 37:30]
  wire  _T_1264 = 8'h3 == _T_1261; // @[Conditional.scala 37:30]
  wire  _GEN_111 = _T_1262 ? regs[55] : _T_1264; // @[Conditional.scala 40:58]
  wire [1:0] _T_1273 = regs[39] + regs[40]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_849 = {{1'd0}, regs[41]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1274 = _T_1273 + _GEN_849; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_850 = {{2'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1275 = _T_1274 + _GEN_850; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_851 = {{3'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1276 = _T_1275 + _GEN_851; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_852 = {{4'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1277 = _T_1276 + _GEN_852; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_853 = {{5'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1278 = _T_1277 + _GEN_853; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_854 = {{6'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1279 = _T_1278 + _GEN_854; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1280 = 8'h2 == _T_1279; // @[Conditional.scala 37:30]
  wire  _T_1282 = 8'h3 == _T_1279; // @[Conditional.scala 37:30]
  wire  _GEN_113 = _T_1280 ? regs[56] : _T_1282; // @[Conditional.scala 40:58]
  wire [1:0] _T_1291 = regs[40] + regs[41]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_855 = {{1'd0}, regs[42]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1292 = _T_1291 + _GEN_855; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_856 = {{2'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1293 = _T_1292 + _GEN_856; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_857 = {{3'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1294 = _T_1293 + _GEN_857; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_858 = {{4'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1295 = _T_1294 + _GEN_858; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_859 = {{5'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1296 = _T_1295 + _GEN_859; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_860 = {{6'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1297 = _T_1296 + _GEN_860; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1298 = 8'h2 == _T_1297; // @[Conditional.scala 37:30]
  wire  _T_1300 = 8'h3 == _T_1297; // @[Conditional.scala 37:30]
  wire  _GEN_115 = _T_1298 ? regs[57] : _T_1300; // @[Conditional.scala 40:58]
  wire [1:0] _T_1309 = regs[41] + regs[42]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_861 = {{1'd0}, regs[43]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1310 = _T_1309 + _GEN_861; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_862 = {{2'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1311 = _T_1310 + _GEN_862; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_863 = {{3'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1312 = _T_1311 + _GEN_863; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_864 = {{4'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1313 = _T_1312 + _GEN_864; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_865 = {{5'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1314 = _T_1313 + _GEN_865; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_866 = {{6'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1315 = _T_1314 + _GEN_866; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1316 = 8'h2 == _T_1315; // @[Conditional.scala 37:30]
  wire  _T_1318 = 8'h3 == _T_1315; // @[Conditional.scala 37:30]
  wire  _GEN_117 = _T_1316 ? regs[58] : _T_1318; // @[Conditional.scala 40:58]
  wire [1:0] _T_1327 = regs[42] + regs[43]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_867 = {{1'd0}, regs[44]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1328 = _T_1327 + _GEN_867; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_868 = {{2'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1329 = _T_1328 + _GEN_868; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_869 = {{3'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1330 = _T_1329 + _GEN_869; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_870 = {{4'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1331 = _T_1330 + _GEN_870; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_871 = {{5'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1332 = _T_1331 + _GEN_871; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_872 = {{6'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1333 = _T_1332 + _GEN_872; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1334 = 8'h2 == _T_1333; // @[Conditional.scala 37:30]
  wire  _T_1336 = 8'h3 == _T_1333; // @[Conditional.scala 37:30]
  wire  _GEN_119 = _T_1334 ? regs[59] : _T_1336; // @[Conditional.scala 40:58]
  wire [1:0] _T_1345 = regs[43] + regs[44]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_873 = {{1'd0}, regs[45]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1346 = _T_1345 + _GEN_873; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_874 = {{2'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1347 = _T_1346 + _GEN_874; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_875 = {{3'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1348 = _T_1347 + _GEN_875; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_876 = {{4'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1349 = _T_1348 + _GEN_876; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_877 = {{5'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1350 = _T_1349 + _GEN_877; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_878 = {{6'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1351 = _T_1350 + _GEN_878; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1352 = 8'h2 == _T_1351; // @[Conditional.scala 37:30]
  wire  _T_1354 = 8'h3 == _T_1351; // @[Conditional.scala 37:30]
  wire  _GEN_121 = _T_1352 ? regs[60] : _T_1354; // @[Conditional.scala 40:58]
  wire [1:0] _T_1363 = regs[44] + regs[45]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_879 = {{1'd0}, regs[46]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1364 = _T_1363 + _GEN_879; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_880 = {{2'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1365 = _T_1364 + _GEN_880; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_881 = {{3'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1366 = _T_1365 + _GEN_881; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_882 = {{4'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1367 = _T_1366 + _GEN_882; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_883 = {{5'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1368 = _T_1367 + _GEN_883; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_884 = {{6'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1369 = _T_1368 + _GEN_884; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1370 = 8'h2 == _T_1369; // @[Conditional.scala 37:30]
  wire  _T_1372 = 8'h3 == _T_1369; // @[Conditional.scala 37:30]
  wire  _GEN_123 = _T_1370 ? regs[61] : _T_1372; // @[Conditional.scala 40:58]
  wire [1:0] _T_1381 = regs[45] + regs[46]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_885 = {{1'd0}, regs[47]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1382 = _T_1381 + _GEN_885; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_886 = {{2'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1383 = _T_1382 + _GEN_886; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_887 = {{3'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1384 = _T_1383 + _GEN_887; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_888 = {{4'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1385 = _T_1384 + _GEN_888; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_889 = {{5'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1386 = _T_1385 + _GEN_889; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_890 = {{6'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1387 = _T_1386 + _GEN_890; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1388 = 8'h2 == _T_1387; // @[Conditional.scala 37:30]
  wire  _T_1390 = 8'h3 == _T_1387; // @[Conditional.scala 37:30]
  wire  _GEN_125 = _T_1388 ? regs[62] : _T_1390; // @[Conditional.scala 40:58]
  wire [1:0] _T_1399 = regs[46] + regs[47]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_891 = {{1'd0}, regs[32]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1400 = _T_1399 + _GEN_891; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_892 = {{2'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1401 = _T_1400 + _GEN_892; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_893 = {{3'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1402 = _T_1401 + _GEN_893; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_894 = {{4'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1403 = _T_1402 + _GEN_894; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_895 = {{5'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1404 = _T_1403 + _GEN_895; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_896 = {{6'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1405 = _T_1404 + _GEN_896; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1406 = 8'h2 == _T_1405; // @[Conditional.scala 37:30]
  wire  _T_1408 = 8'h3 == _T_1405; // @[Conditional.scala 37:30]
  wire  _GEN_127 = _T_1406 ? regs[63] : _T_1408; // @[Conditional.scala 40:58]
  wire [1:0] _T_1417 = regs[63] + regs[48]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_897 = {{1'd0}, regs[49]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1418 = _T_1417 + _GEN_897; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_898 = {{2'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1419 = _T_1418 + _GEN_898; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_899 = {{3'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1420 = _T_1419 + _GEN_899; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_900 = {{4'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1421 = _T_1420 + _GEN_900; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_901 = {{5'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1422 = _T_1421 + _GEN_901; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_902 = {{6'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1423 = _T_1422 + _GEN_902; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1424 = 8'h2 == _T_1423; // @[Conditional.scala 37:30]
  wire  _T_1426 = 8'h3 == _T_1423; // @[Conditional.scala 37:30]
  wire  _GEN_129 = _T_1424 ? regs[64] : _T_1426; // @[Conditional.scala 40:58]
  wire [1:0] _T_1435 = regs[48] + regs[49]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_903 = {{1'd0}, regs[50]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1436 = _T_1435 + _GEN_903; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_904 = {{2'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1437 = _T_1436 + _GEN_904; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_905 = {{3'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1438 = _T_1437 + _GEN_905; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_906 = {{4'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1439 = _T_1438 + _GEN_906; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_907 = {{5'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1440 = _T_1439 + _GEN_907; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_908 = {{6'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1441 = _T_1440 + _GEN_908; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1442 = 8'h2 == _T_1441; // @[Conditional.scala 37:30]
  wire  _T_1444 = 8'h3 == _T_1441; // @[Conditional.scala 37:30]
  wire  _GEN_131 = _T_1442 ? regs[65] : _T_1444; // @[Conditional.scala 40:58]
  wire [1:0] _T_1453 = regs[49] + regs[50]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_909 = {{1'd0}, regs[51]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1454 = _T_1453 + _GEN_909; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_910 = {{2'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1455 = _T_1454 + _GEN_910; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_911 = {{3'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1456 = _T_1455 + _GEN_911; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_912 = {{4'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1457 = _T_1456 + _GEN_912; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_913 = {{5'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1458 = _T_1457 + _GEN_913; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_914 = {{6'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1459 = _T_1458 + _GEN_914; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1460 = 8'h2 == _T_1459; // @[Conditional.scala 37:30]
  wire  _T_1462 = 8'h3 == _T_1459; // @[Conditional.scala 37:30]
  wire  _GEN_133 = _T_1460 ? regs[66] : _T_1462; // @[Conditional.scala 40:58]
  wire [1:0] _T_1471 = regs[50] + regs[51]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_915 = {{1'd0}, regs[52]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1472 = _T_1471 + _GEN_915; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_916 = {{2'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1473 = _T_1472 + _GEN_916; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_917 = {{3'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1474 = _T_1473 + _GEN_917; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_918 = {{4'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1475 = _T_1474 + _GEN_918; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_919 = {{5'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1476 = _T_1475 + _GEN_919; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_920 = {{6'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1477 = _T_1476 + _GEN_920; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1478 = 8'h2 == _T_1477; // @[Conditional.scala 37:30]
  wire  _T_1480 = 8'h3 == _T_1477; // @[Conditional.scala 37:30]
  wire  _GEN_135 = _T_1478 ? regs[67] : _T_1480; // @[Conditional.scala 40:58]
  wire [1:0] _T_1489 = regs[51] + regs[52]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_921 = {{1'd0}, regs[53]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1490 = _T_1489 + _GEN_921; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_922 = {{2'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1491 = _T_1490 + _GEN_922; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_923 = {{3'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1492 = _T_1491 + _GEN_923; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_924 = {{4'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1493 = _T_1492 + _GEN_924; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_925 = {{5'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1494 = _T_1493 + _GEN_925; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_926 = {{6'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1495 = _T_1494 + _GEN_926; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1496 = 8'h2 == _T_1495; // @[Conditional.scala 37:30]
  wire  _T_1498 = 8'h3 == _T_1495; // @[Conditional.scala 37:30]
  wire  _GEN_137 = _T_1496 ? regs[68] : _T_1498; // @[Conditional.scala 40:58]
  wire [1:0] _T_1507 = regs[52] + regs[53]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_927 = {{1'd0}, regs[54]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1508 = _T_1507 + _GEN_927; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_928 = {{2'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1509 = _T_1508 + _GEN_928; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_929 = {{3'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1510 = _T_1509 + _GEN_929; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_930 = {{4'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1511 = _T_1510 + _GEN_930; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_931 = {{5'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1512 = _T_1511 + _GEN_931; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_932 = {{6'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1513 = _T_1512 + _GEN_932; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1514 = 8'h2 == _T_1513; // @[Conditional.scala 37:30]
  wire  _T_1516 = 8'h3 == _T_1513; // @[Conditional.scala 37:30]
  wire  _GEN_139 = _T_1514 ? regs[69] : _T_1516; // @[Conditional.scala 40:58]
  wire [1:0] _T_1525 = regs[53] + regs[54]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_933 = {{1'd0}, regs[55]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1526 = _T_1525 + _GEN_933; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_934 = {{2'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1527 = _T_1526 + _GEN_934; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_935 = {{3'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1528 = _T_1527 + _GEN_935; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_936 = {{4'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1529 = _T_1528 + _GEN_936; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_937 = {{5'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1530 = _T_1529 + _GEN_937; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_938 = {{6'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1531 = _T_1530 + _GEN_938; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1532 = 8'h2 == _T_1531; // @[Conditional.scala 37:30]
  wire  _T_1534 = 8'h3 == _T_1531; // @[Conditional.scala 37:30]
  wire  _GEN_141 = _T_1532 ? regs[70] : _T_1534; // @[Conditional.scala 40:58]
  wire [1:0] _T_1543 = regs[54] + regs[55]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_939 = {{1'd0}, regs[56]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1544 = _T_1543 + _GEN_939; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_940 = {{2'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1545 = _T_1544 + _GEN_940; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_941 = {{3'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1546 = _T_1545 + _GEN_941; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_942 = {{4'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1547 = _T_1546 + _GEN_942; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_943 = {{5'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1548 = _T_1547 + _GEN_943; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_944 = {{6'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1549 = _T_1548 + _GEN_944; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1550 = 8'h2 == _T_1549; // @[Conditional.scala 37:30]
  wire  _T_1552 = 8'h3 == _T_1549; // @[Conditional.scala 37:30]
  wire  _GEN_143 = _T_1550 ? regs[71] : _T_1552; // @[Conditional.scala 40:58]
  wire [1:0] _T_1561 = regs[55] + regs[56]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_945 = {{1'd0}, regs[57]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1562 = _T_1561 + _GEN_945; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_946 = {{2'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1563 = _T_1562 + _GEN_946; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_947 = {{3'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1564 = _T_1563 + _GEN_947; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_948 = {{4'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1565 = _T_1564 + _GEN_948; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_949 = {{5'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1566 = _T_1565 + _GEN_949; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_950 = {{6'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1567 = _T_1566 + _GEN_950; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1568 = 8'h2 == _T_1567; // @[Conditional.scala 37:30]
  wire  _T_1570 = 8'h3 == _T_1567; // @[Conditional.scala 37:30]
  wire  _GEN_145 = _T_1568 ? regs[72] : _T_1570; // @[Conditional.scala 40:58]
  wire [1:0] _T_1579 = regs[56] + regs[57]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_951 = {{1'd0}, regs[58]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1580 = _T_1579 + _GEN_951; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_952 = {{2'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1581 = _T_1580 + _GEN_952; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_953 = {{3'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1582 = _T_1581 + _GEN_953; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_954 = {{4'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1583 = _T_1582 + _GEN_954; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_955 = {{5'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1584 = _T_1583 + _GEN_955; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_956 = {{6'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1585 = _T_1584 + _GEN_956; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1586 = 8'h2 == _T_1585; // @[Conditional.scala 37:30]
  wire  _T_1588 = 8'h3 == _T_1585; // @[Conditional.scala 37:30]
  wire  _GEN_147 = _T_1586 ? regs[73] : _T_1588; // @[Conditional.scala 40:58]
  wire [1:0] _T_1597 = regs[57] + regs[58]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_957 = {{1'd0}, regs[59]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1598 = _T_1597 + _GEN_957; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_958 = {{2'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1599 = _T_1598 + _GEN_958; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_959 = {{3'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1600 = _T_1599 + _GEN_959; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_960 = {{4'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1601 = _T_1600 + _GEN_960; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_961 = {{5'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1602 = _T_1601 + _GEN_961; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_962 = {{6'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1603 = _T_1602 + _GEN_962; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1604 = 8'h2 == _T_1603; // @[Conditional.scala 37:30]
  wire  _T_1606 = 8'h3 == _T_1603; // @[Conditional.scala 37:30]
  wire  _GEN_149 = _T_1604 ? regs[74] : _T_1606; // @[Conditional.scala 40:58]
  wire [1:0] _T_1615 = regs[58] + regs[59]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_963 = {{1'd0}, regs[60]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1616 = _T_1615 + _GEN_963; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_964 = {{2'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1617 = _T_1616 + _GEN_964; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_965 = {{3'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1618 = _T_1617 + _GEN_965; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_966 = {{4'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1619 = _T_1618 + _GEN_966; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_967 = {{5'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1620 = _T_1619 + _GEN_967; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_968 = {{6'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1621 = _T_1620 + _GEN_968; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1622 = 8'h2 == _T_1621; // @[Conditional.scala 37:30]
  wire  _T_1624 = 8'h3 == _T_1621; // @[Conditional.scala 37:30]
  wire  _GEN_151 = _T_1622 ? regs[75] : _T_1624; // @[Conditional.scala 40:58]
  wire [1:0] _T_1633 = regs[59] + regs[60]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_969 = {{1'd0}, regs[61]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1634 = _T_1633 + _GEN_969; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_970 = {{2'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1635 = _T_1634 + _GEN_970; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_971 = {{3'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1636 = _T_1635 + _GEN_971; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_972 = {{4'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1637 = _T_1636 + _GEN_972; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_973 = {{5'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1638 = _T_1637 + _GEN_973; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_974 = {{6'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1639 = _T_1638 + _GEN_974; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1640 = 8'h2 == _T_1639; // @[Conditional.scala 37:30]
  wire  _T_1642 = 8'h3 == _T_1639; // @[Conditional.scala 37:30]
  wire  _GEN_153 = _T_1640 ? regs[76] : _T_1642; // @[Conditional.scala 40:58]
  wire [1:0] _T_1651 = regs[60] + regs[61]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_975 = {{1'd0}, regs[62]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1652 = _T_1651 + _GEN_975; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_976 = {{2'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1653 = _T_1652 + _GEN_976; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_977 = {{3'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1654 = _T_1653 + _GEN_977; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_978 = {{4'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1655 = _T_1654 + _GEN_978; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_979 = {{5'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1656 = _T_1655 + _GEN_979; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_980 = {{6'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1657 = _T_1656 + _GEN_980; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1658 = 8'h2 == _T_1657; // @[Conditional.scala 37:30]
  wire  _T_1660 = 8'h3 == _T_1657; // @[Conditional.scala 37:30]
  wire  _GEN_155 = _T_1658 ? regs[77] : _T_1660; // @[Conditional.scala 40:58]
  wire [1:0] _T_1669 = regs[61] + regs[62]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_981 = {{1'd0}, regs[63]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1670 = _T_1669 + _GEN_981; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_982 = {{2'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1671 = _T_1670 + _GEN_982; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_983 = {{3'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1672 = _T_1671 + _GEN_983; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_984 = {{4'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1673 = _T_1672 + _GEN_984; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_985 = {{5'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1674 = _T_1673 + _GEN_985; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_986 = {{6'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1675 = _T_1674 + _GEN_986; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1676 = 8'h2 == _T_1675; // @[Conditional.scala 37:30]
  wire  _T_1678 = 8'h3 == _T_1675; // @[Conditional.scala 37:30]
  wire  _GEN_157 = _T_1676 ? regs[78] : _T_1678; // @[Conditional.scala 40:58]
  wire [1:0] _T_1687 = regs[62] + regs[63]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_987 = {{1'd0}, regs[48]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1688 = _T_1687 + _GEN_987; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_988 = {{2'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1689 = _T_1688 + _GEN_988; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_989 = {{3'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1690 = _T_1689 + _GEN_989; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_990 = {{4'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1691 = _T_1690 + _GEN_990; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_991 = {{5'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1692 = _T_1691 + _GEN_991; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_992 = {{6'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1693 = _T_1692 + _GEN_992; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1694 = 8'h2 == _T_1693; // @[Conditional.scala 37:30]
  wire  _T_1696 = 8'h3 == _T_1693; // @[Conditional.scala 37:30]
  wire  _GEN_159 = _T_1694 ? regs[79] : _T_1696; // @[Conditional.scala 40:58]
  wire [1:0] _T_1705 = regs[79] + regs[64]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_993 = {{1'd0}, regs[65]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1706 = _T_1705 + _GEN_993; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_994 = {{2'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1707 = _T_1706 + _GEN_994; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_995 = {{3'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1708 = _T_1707 + _GEN_995; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_996 = {{4'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1709 = _T_1708 + _GEN_996; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_997 = {{5'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1710 = _T_1709 + _GEN_997; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_998 = {{6'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1711 = _T_1710 + _GEN_998; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1712 = 8'h2 == _T_1711; // @[Conditional.scala 37:30]
  wire  _T_1714 = 8'h3 == _T_1711; // @[Conditional.scala 37:30]
  wire  _GEN_161 = _T_1712 ? regs[80] : _T_1714; // @[Conditional.scala 40:58]
  wire [1:0] _T_1723 = regs[64] + regs[65]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_999 = {{1'd0}, regs[66]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1724 = _T_1723 + _GEN_999; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1000 = {{2'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1725 = _T_1724 + _GEN_1000; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1001 = {{3'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1726 = _T_1725 + _GEN_1001; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1002 = {{4'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1727 = _T_1726 + _GEN_1002; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1003 = {{5'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1728 = _T_1727 + _GEN_1003; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1004 = {{6'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1729 = _T_1728 + _GEN_1004; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1730 = 8'h2 == _T_1729; // @[Conditional.scala 37:30]
  wire  _T_1732 = 8'h3 == _T_1729; // @[Conditional.scala 37:30]
  wire  _GEN_163 = _T_1730 ? regs[81] : _T_1732; // @[Conditional.scala 40:58]
  wire [1:0] _T_1741 = regs[65] + regs[66]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1005 = {{1'd0}, regs[67]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1742 = _T_1741 + _GEN_1005; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1006 = {{2'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1743 = _T_1742 + _GEN_1006; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1007 = {{3'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1744 = _T_1743 + _GEN_1007; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1008 = {{4'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1745 = _T_1744 + _GEN_1008; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1009 = {{5'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1746 = _T_1745 + _GEN_1009; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1010 = {{6'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1747 = _T_1746 + _GEN_1010; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1748 = 8'h2 == _T_1747; // @[Conditional.scala 37:30]
  wire  _T_1750 = 8'h3 == _T_1747; // @[Conditional.scala 37:30]
  wire  _GEN_165 = _T_1748 ? regs[82] : _T_1750; // @[Conditional.scala 40:58]
  wire [1:0] _T_1759 = regs[66] + regs[67]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1011 = {{1'd0}, regs[68]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1760 = _T_1759 + _GEN_1011; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1012 = {{2'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1761 = _T_1760 + _GEN_1012; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1013 = {{3'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1762 = _T_1761 + _GEN_1013; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1014 = {{4'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1763 = _T_1762 + _GEN_1014; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1015 = {{5'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1764 = _T_1763 + _GEN_1015; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1016 = {{6'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1765 = _T_1764 + _GEN_1016; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1766 = 8'h2 == _T_1765; // @[Conditional.scala 37:30]
  wire  _T_1768 = 8'h3 == _T_1765; // @[Conditional.scala 37:30]
  wire  _GEN_167 = _T_1766 ? regs[83] : _T_1768; // @[Conditional.scala 40:58]
  wire [1:0] _T_1777 = regs[67] + regs[68]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1017 = {{1'd0}, regs[69]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1778 = _T_1777 + _GEN_1017; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1018 = {{2'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1779 = _T_1778 + _GEN_1018; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1019 = {{3'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1780 = _T_1779 + _GEN_1019; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1020 = {{4'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1781 = _T_1780 + _GEN_1020; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1021 = {{5'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1782 = _T_1781 + _GEN_1021; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1022 = {{6'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1783 = _T_1782 + _GEN_1022; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1784 = 8'h2 == _T_1783; // @[Conditional.scala 37:30]
  wire  _T_1786 = 8'h3 == _T_1783; // @[Conditional.scala 37:30]
  wire  _GEN_169 = _T_1784 ? regs[84] : _T_1786; // @[Conditional.scala 40:58]
  wire [1:0] _T_1795 = regs[68] + regs[69]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1023 = {{1'd0}, regs[70]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1796 = _T_1795 + _GEN_1023; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1024 = {{2'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1797 = _T_1796 + _GEN_1024; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1025 = {{3'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1798 = _T_1797 + _GEN_1025; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1026 = {{4'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1799 = _T_1798 + _GEN_1026; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1027 = {{5'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1800 = _T_1799 + _GEN_1027; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1028 = {{6'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1801 = _T_1800 + _GEN_1028; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1802 = 8'h2 == _T_1801; // @[Conditional.scala 37:30]
  wire  _T_1804 = 8'h3 == _T_1801; // @[Conditional.scala 37:30]
  wire  _GEN_171 = _T_1802 ? regs[85] : _T_1804; // @[Conditional.scala 40:58]
  wire [1:0] _T_1813 = regs[69] + regs[70]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1029 = {{1'd0}, regs[71]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1814 = _T_1813 + _GEN_1029; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1030 = {{2'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1815 = _T_1814 + _GEN_1030; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1031 = {{3'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1816 = _T_1815 + _GEN_1031; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1032 = {{4'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1817 = _T_1816 + _GEN_1032; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1033 = {{5'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1818 = _T_1817 + _GEN_1033; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1034 = {{6'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1819 = _T_1818 + _GEN_1034; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1820 = 8'h2 == _T_1819; // @[Conditional.scala 37:30]
  wire  _T_1822 = 8'h3 == _T_1819; // @[Conditional.scala 37:30]
  wire  _GEN_173 = _T_1820 ? regs[86] : _T_1822; // @[Conditional.scala 40:58]
  wire [1:0] _T_1831 = regs[70] + regs[71]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1035 = {{1'd0}, regs[72]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1832 = _T_1831 + _GEN_1035; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1036 = {{2'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1833 = _T_1832 + _GEN_1036; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1037 = {{3'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1834 = _T_1833 + _GEN_1037; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1038 = {{4'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1835 = _T_1834 + _GEN_1038; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1039 = {{5'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1836 = _T_1835 + _GEN_1039; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1040 = {{6'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1837 = _T_1836 + _GEN_1040; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1838 = 8'h2 == _T_1837; // @[Conditional.scala 37:30]
  wire  _T_1840 = 8'h3 == _T_1837; // @[Conditional.scala 37:30]
  wire  _GEN_175 = _T_1838 ? regs[87] : _T_1840; // @[Conditional.scala 40:58]
  wire [1:0] _T_1849 = regs[71] + regs[72]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1041 = {{1'd0}, regs[73]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1850 = _T_1849 + _GEN_1041; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1042 = {{2'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1851 = _T_1850 + _GEN_1042; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1043 = {{3'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1852 = _T_1851 + _GEN_1043; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1044 = {{4'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1853 = _T_1852 + _GEN_1044; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1045 = {{5'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1854 = _T_1853 + _GEN_1045; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1046 = {{6'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1855 = _T_1854 + _GEN_1046; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1856 = 8'h2 == _T_1855; // @[Conditional.scala 37:30]
  wire  _T_1858 = 8'h3 == _T_1855; // @[Conditional.scala 37:30]
  wire  _GEN_177 = _T_1856 ? regs[88] : _T_1858; // @[Conditional.scala 40:58]
  wire [1:0] _T_1867 = regs[72] + regs[73]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1047 = {{1'd0}, regs[74]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1868 = _T_1867 + _GEN_1047; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1048 = {{2'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1869 = _T_1868 + _GEN_1048; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1049 = {{3'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1870 = _T_1869 + _GEN_1049; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1050 = {{4'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1871 = _T_1870 + _GEN_1050; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1051 = {{5'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1872 = _T_1871 + _GEN_1051; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1052 = {{6'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1873 = _T_1872 + _GEN_1052; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1874 = 8'h2 == _T_1873; // @[Conditional.scala 37:30]
  wire  _T_1876 = 8'h3 == _T_1873; // @[Conditional.scala 37:30]
  wire  _GEN_179 = _T_1874 ? regs[89] : _T_1876; // @[Conditional.scala 40:58]
  wire [1:0] _T_1885 = regs[73] + regs[74]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1053 = {{1'd0}, regs[75]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1886 = _T_1885 + _GEN_1053; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1054 = {{2'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1887 = _T_1886 + _GEN_1054; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1055 = {{3'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1888 = _T_1887 + _GEN_1055; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1056 = {{4'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1889 = _T_1888 + _GEN_1056; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1057 = {{5'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1890 = _T_1889 + _GEN_1057; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1058 = {{6'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1891 = _T_1890 + _GEN_1058; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1892 = 8'h2 == _T_1891; // @[Conditional.scala 37:30]
  wire  _T_1894 = 8'h3 == _T_1891; // @[Conditional.scala 37:30]
  wire  _GEN_181 = _T_1892 ? regs[90] : _T_1894; // @[Conditional.scala 40:58]
  wire [1:0] _T_1903 = regs[74] + regs[75]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1059 = {{1'd0}, regs[76]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1904 = _T_1903 + _GEN_1059; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1060 = {{2'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1905 = _T_1904 + _GEN_1060; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1061 = {{3'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1906 = _T_1905 + _GEN_1061; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1062 = {{4'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1907 = _T_1906 + _GEN_1062; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1063 = {{5'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1908 = _T_1907 + _GEN_1063; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1064 = {{6'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1909 = _T_1908 + _GEN_1064; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1910 = 8'h2 == _T_1909; // @[Conditional.scala 37:30]
  wire  _T_1912 = 8'h3 == _T_1909; // @[Conditional.scala 37:30]
  wire  _GEN_183 = _T_1910 ? regs[91] : _T_1912; // @[Conditional.scala 40:58]
  wire [1:0] _T_1921 = regs[75] + regs[76]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1065 = {{1'd0}, regs[77]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1922 = _T_1921 + _GEN_1065; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1066 = {{2'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1923 = _T_1922 + _GEN_1066; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1067 = {{3'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1924 = _T_1923 + _GEN_1067; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1068 = {{4'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1925 = _T_1924 + _GEN_1068; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1069 = {{5'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1926 = _T_1925 + _GEN_1069; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1070 = {{6'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1927 = _T_1926 + _GEN_1070; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1928 = 8'h2 == _T_1927; // @[Conditional.scala 37:30]
  wire  _T_1930 = 8'h3 == _T_1927; // @[Conditional.scala 37:30]
  wire  _GEN_185 = _T_1928 ? regs[92] : _T_1930; // @[Conditional.scala 40:58]
  wire [1:0] _T_1939 = regs[76] + regs[77]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1071 = {{1'd0}, regs[78]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1940 = _T_1939 + _GEN_1071; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1072 = {{2'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1941 = _T_1940 + _GEN_1072; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1073 = {{3'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1942 = _T_1941 + _GEN_1073; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1074 = {{4'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1943 = _T_1942 + _GEN_1074; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1075 = {{5'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1944 = _T_1943 + _GEN_1075; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1076 = {{6'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1945 = _T_1944 + _GEN_1076; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1946 = 8'h2 == _T_1945; // @[Conditional.scala 37:30]
  wire  _T_1948 = 8'h3 == _T_1945; // @[Conditional.scala 37:30]
  wire  _GEN_187 = _T_1946 ? regs[93] : _T_1948; // @[Conditional.scala 40:58]
  wire [1:0] _T_1957 = regs[77] + regs[78]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1077 = {{1'd0}, regs[79]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1958 = _T_1957 + _GEN_1077; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1078 = {{2'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1959 = _T_1958 + _GEN_1078; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1079 = {{3'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1960 = _T_1959 + _GEN_1079; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1080 = {{4'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1961 = _T_1960 + _GEN_1080; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1081 = {{5'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1962 = _T_1961 + _GEN_1081; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1082 = {{6'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1963 = _T_1962 + _GEN_1082; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1964 = 8'h2 == _T_1963; // @[Conditional.scala 37:30]
  wire  _T_1966 = 8'h3 == _T_1963; // @[Conditional.scala 37:30]
  wire  _GEN_189 = _T_1964 ? regs[94] : _T_1966; // @[Conditional.scala 40:58]
  wire [1:0] _T_1975 = regs[78] + regs[79]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1083 = {{1'd0}, regs[64]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1976 = _T_1975 + _GEN_1083; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1084 = {{2'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1977 = _T_1976 + _GEN_1084; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1085 = {{3'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1978 = _T_1977 + _GEN_1085; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1086 = {{4'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1979 = _T_1978 + _GEN_1086; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1087 = {{5'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1980 = _T_1979 + _GEN_1087; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1088 = {{6'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1981 = _T_1980 + _GEN_1088; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_1982 = 8'h2 == _T_1981; // @[Conditional.scala 37:30]
  wire  _T_1984 = 8'h3 == _T_1981; // @[Conditional.scala 37:30]
  wire  _GEN_191 = _T_1982 ? regs[95] : _T_1984; // @[Conditional.scala 40:58]
  wire [1:0] _T_1993 = regs[95] + regs[80]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1089 = {{1'd0}, regs[81]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_1994 = _T_1993 + _GEN_1089; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1090 = {{2'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_1995 = _T_1994 + _GEN_1090; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1091 = {{3'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_1996 = _T_1995 + _GEN_1091; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1092 = {{4'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_1997 = _T_1996 + _GEN_1092; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1093 = {{5'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_1998 = _T_1997 + _GEN_1093; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1094 = {{6'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_1999 = _T_1998 + _GEN_1094; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2000 = 8'h2 == _T_1999; // @[Conditional.scala 37:30]
  wire  _T_2002 = 8'h3 == _T_1999; // @[Conditional.scala 37:30]
  wire  _GEN_193 = _T_2000 ? regs[96] : _T_2002; // @[Conditional.scala 40:58]
  wire [1:0] _T_2011 = regs[80] + regs[81]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1095 = {{1'd0}, regs[82]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2012 = _T_2011 + _GEN_1095; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1096 = {{2'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2013 = _T_2012 + _GEN_1096; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1097 = {{3'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2014 = _T_2013 + _GEN_1097; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1098 = {{4'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2015 = _T_2014 + _GEN_1098; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1099 = {{5'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2016 = _T_2015 + _GEN_1099; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1100 = {{6'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2017 = _T_2016 + _GEN_1100; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2018 = 8'h2 == _T_2017; // @[Conditional.scala 37:30]
  wire  _T_2020 = 8'h3 == _T_2017; // @[Conditional.scala 37:30]
  wire  _GEN_195 = _T_2018 ? regs[97] : _T_2020; // @[Conditional.scala 40:58]
  wire [1:0] _T_2029 = regs[81] + regs[82]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1101 = {{1'd0}, regs[83]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2030 = _T_2029 + _GEN_1101; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1102 = {{2'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2031 = _T_2030 + _GEN_1102; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1103 = {{3'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2032 = _T_2031 + _GEN_1103; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1104 = {{4'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2033 = _T_2032 + _GEN_1104; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1105 = {{5'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2034 = _T_2033 + _GEN_1105; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1106 = {{6'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2035 = _T_2034 + _GEN_1106; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2036 = 8'h2 == _T_2035; // @[Conditional.scala 37:30]
  wire  _T_2038 = 8'h3 == _T_2035; // @[Conditional.scala 37:30]
  wire  _GEN_197 = _T_2036 ? regs[98] : _T_2038; // @[Conditional.scala 40:58]
  wire [1:0] _T_2047 = regs[82] + regs[83]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1107 = {{1'd0}, regs[84]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2048 = _T_2047 + _GEN_1107; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1108 = {{2'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2049 = _T_2048 + _GEN_1108; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1109 = {{3'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2050 = _T_2049 + _GEN_1109; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1110 = {{4'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2051 = _T_2050 + _GEN_1110; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1111 = {{5'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2052 = _T_2051 + _GEN_1111; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1112 = {{6'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2053 = _T_2052 + _GEN_1112; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2054 = 8'h2 == _T_2053; // @[Conditional.scala 37:30]
  wire  _T_2056 = 8'h3 == _T_2053; // @[Conditional.scala 37:30]
  wire  _GEN_199 = _T_2054 ? regs[99] : _T_2056; // @[Conditional.scala 40:58]
  wire [1:0] _T_2065 = regs[83] + regs[84]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1113 = {{1'd0}, regs[85]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2066 = _T_2065 + _GEN_1113; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1114 = {{2'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2067 = _T_2066 + _GEN_1114; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1115 = {{3'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2068 = _T_2067 + _GEN_1115; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1116 = {{4'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2069 = _T_2068 + _GEN_1116; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1117 = {{5'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2070 = _T_2069 + _GEN_1117; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1118 = {{6'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2071 = _T_2070 + _GEN_1118; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2072 = 8'h2 == _T_2071; // @[Conditional.scala 37:30]
  wire  _T_2074 = 8'h3 == _T_2071; // @[Conditional.scala 37:30]
  wire  _GEN_201 = _T_2072 ? regs[100] : _T_2074; // @[Conditional.scala 40:58]
  wire [1:0] _T_2083 = regs[84] + regs[85]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1119 = {{1'd0}, regs[86]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2084 = _T_2083 + _GEN_1119; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1120 = {{2'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2085 = _T_2084 + _GEN_1120; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1121 = {{3'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2086 = _T_2085 + _GEN_1121; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1122 = {{4'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2087 = _T_2086 + _GEN_1122; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1123 = {{5'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2088 = _T_2087 + _GEN_1123; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1124 = {{6'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2089 = _T_2088 + _GEN_1124; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2090 = 8'h2 == _T_2089; // @[Conditional.scala 37:30]
  wire  _T_2092 = 8'h3 == _T_2089; // @[Conditional.scala 37:30]
  wire  _GEN_203 = _T_2090 ? regs[101] : _T_2092; // @[Conditional.scala 40:58]
  wire [1:0] _T_2101 = regs[85] + regs[86]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1125 = {{1'd0}, regs[87]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2102 = _T_2101 + _GEN_1125; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1126 = {{2'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2103 = _T_2102 + _GEN_1126; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1127 = {{3'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2104 = _T_2103 + _GEN_1127; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1128 = {{4'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2105 = _T_2104 + _GEN_1128; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1129 = {{5'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2106 = _T_2105 + _GEN_1129; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1130 = {{6'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2107 = _T_2106 + _GEN_1130; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2108 = 8'h2 == _T_2107; // @[Conditional.scala 37:30]
  wire  _T_2110 = 8'h3 == _T_2107; // @[Conditional.scala 37:30]
  wire  _GEN_205 = _T_2108 ? regs[102] : _T_2110; // @[Conditional.scala 40:58]
  wire [1:0] _T_2119 = regs[86] + regs[87]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1131 = {{1'd0}, regs[88]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2120 = _T_2119 + _GEN_1131; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1132 = {{2'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2121 = _T_2120 + _GEN_1132; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1133 = {{3'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2122 = _T_2121 + _GEN_1133; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1134 = {{4'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2123 = _T_2122 + _GEN_1134; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1135 = {{5'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2124 = _T_2123 + _GEN_1135; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1136 = {{6'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2125 = _T_2124 + _GEN_1136; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2126 = 8'h2 == _T_2125; // @[Conditional.scala 37:30]
  wire  _T_2128 = 8'h3 == _T_2125; // @[Conditional.scala 37:30]
  wire  _GEN_207 = _T_2126 ? regs[103] : _T_2128; // @[Conditional.scala 40:58]
  wire [1:0] _T_2137 = regs[87] + regs[88]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1137 = {{1'd0}, regs[89]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2138 = _T_2137 + _GEN_1137; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1138 = {{2'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2139 = _T_2138 + _GEN_1138; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1139 = {{3'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2140 = _T_2139 + _GEN_1139; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1140 = {{4'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2141 = _T_2140 + _GEN_1140; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1141 = {{5'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2142 = _T_2141 + _GEN_1141; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1142 = {{6'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2143 = _T_2142 + _GEN_1142; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2144 = 8'h2 == _T_2143; // @[Conditional.scala 37:30]
  wire  _T_2146 = 8'h3 == _T_2143; // @[Conditional.scala 37:30]
  wire  _GEN_209 = _T_2144 ? regs[104] : _T_2146; // @[Conditional.scala 40:58]
  wire [1:0] _T_2155 = regs[88] + regs[89]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1143 = {{1'd0}, regs[90]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2156 = _T_2155 + _GEN_1143; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1144 = {{2'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2157 = _T_2156 + _GEN_1144; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1145 = {{3'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2158 = _T_2157 + _GEN_1145; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1146 = {{4'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2159 = _T_2158 + _GEN_1146; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1147 = {{5'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2160 = _T_2159 + _GEN_1147; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1148 = {{6'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2161 = _T_2160 + _GEN_1148; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2162 = 8'h2 == _T_2161; // @[Conditional.scala 37:30]
  wire  _T_2164 = 8'h3 == _T_2161; // @[Conditional.scala 37:30]
  wire  _GEN_211 = _T_2162 ? regs[105] : _T_2164; // @[Conditional.scala 40:58]
  wire [1:0] _T_2173 = regs[89] + regs[90]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1149 = {{1'd0}, regs[91]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2174 = _T_2173 + _GEN_1149; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1150 = {{2'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2175 = _T_2174 + _GEN_1150; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1151 = {{3'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2176 = _T_2175 + _GEN_1151; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1152 = {{4'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2177 = _T_2176 + _GEN_1152; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1153 = {{5'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2178 = _T_2177 + _GEN_1153; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1154 = {{6'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2179 = _T_2178 + _GEN_1154; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2180 = 8'h2 == _T_2179; // @[Conditional.scala 37:30]
  wire  _T_2182 = 8'h3 == _T_2179; // @[Conditional.scala 37:30]
  wire  _GEN_213 = _T_2180 ? regs[106] : _T_2182; // @[Conditional.scala 40:58]
  wire [1:0] _T_2191 = regs[90] + regs[91]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1155 = {{1'd0}, regs[92]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2192 = _T_2191 + _GEN_1155; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1156 = {{2'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2193 = _T_2192 + _GEN_1156; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1157 = {{3'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2194 = _T_2193 + _GEN_1157; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1158 = {{4'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2195 = _T_2194 + _GEN_1158; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1159 = {{5'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2196 = _T_2195 + _GEN_1159; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1160 = {{6'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2197 = _T_2196 + _GEN_1160; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2198 = 8'h2 == _T_2197; // @[Conditional.scala 37:30]
  wire  _T_2200 = 8'h3 == _T_2197; // @[Conditional.scala 37:30]
  wire  _GEN_215 = _T_2198 ? regs[107] : _T_2200; // @[Conditional.scala 40:58]
  wire [1:0] _T_2209 = regs[91] + regs[92]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1161 = {{1'd0}, regs[93]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2210 = _T_2209 + _GEN_1161; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1162 = {{2'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2211 = _T_2210 + _GEN_1162; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1163 = {{3'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2212 = _T_2211 + _GEN_1163; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1164 = {{4'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2213 = _T_2212 + _GEN_1164; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1165 = {{5'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2214 = _T_2213 + _GEN_1165; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1166 = {{6'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2215 = _T_2214 + _GEN_1166; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2216 = 8'h2 == _T_2215; // @[Conditional.scala 37:30]
  wire  _T_2218 = 8'h3 == _T_2215; // @[Conditional.scala 37:30]
  wire  _GEN_217 = _T_2216 ? regs[108] : _T_2218; // @[Conditional.scala 40:58]
  wire [1:0] _T_2227 = regs[92] + regs[93]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1167 = {{1'd0}, regs[94]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2228 = _T_2227 + _GEN_1167; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1168 = {{2'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2229 = _T_2228 + _GEN_1168; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1169 = {{3'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2230 = _T_2229 + _GEN_1169; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1170 = {{4'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2231 = _T_2230 + _GEN_1170; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1171 = {{5'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2232 = _T_2231 + _GEN_1171; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1172 = {{6'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2233 = _T_2232 + _GEN_1172; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2234 = 8'h2 == _T_2233; // @[Conditional.scala 37:30]
  wire  _T_2236 = 8'h3 == _T_2233; // @[Conditional.scala 37:30]
  wire  _GEN_219 = _T_2234 ? regs[109] : _T_2236; // @[Conditional.scala 40:58]
  wire [1:0] _T_2245 = regs[93] + regs[94]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1173 = {{1'd0}, regs[95]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2246 = _T_2245 + _GEN_1173; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1174 = {{2'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2247 = _T_2246 + _GEN_1174; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1175 = {{3'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2248 = _T_2247 + _GEN_1175; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1176 = {{4'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2249 = _T_2248 + _GEN_1176; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1177 = {{5'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2250 = _T_2249 + _GEN_1177; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1178 = {{6'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2251 = _T_2250 + _GEN_1178; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2252 = 8'h2 == _T_2251; // @[Conditional.scala 37:30]
  wire  _T_2254 = 8'h3 == _T_2251; // @[Conditional.scala 37:30]
  wire  _GEN_221 = _T_2252 ? regs[110] : _T_2254; // @[Conditional.scala 40:58]
  wire [1:0] _T_2263 = regs[94] + regs[95]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1179 = {{1'd0}, regs[80]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2264 = _T_2263 + _GEN_1179; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1180 = {{2'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2265 = _T_2264 + _GEN_1180; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1181 = {{3'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2266 = _T_2265 + _GEN_1181; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1182 = {{4'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2267 = _T_2266 + _GEN_1182; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1183 = {{5'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2268 = _T_2267 + _GEN_1183; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1184 = {{6'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2269 = _T_2268 + _GEN_1184; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2270 = 8'h2 == _T_2269; // @[Conditional.scala 37:30]
  wire  _T_2272 = 8'h3 == _T_2269; // @[Conditional.scala 37:30]
  wire  _GEN_223 = _T_2270 ? regs[111] : _T_2272; // @[Conditional.scala 40:58]
  wire [1:0] _T_2281 = regs[111] + regs[96]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1185 = {{1'd0}, regs[97]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2282 = _T_2281 + _GEN_1185; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1186 = {{2'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2283 = _T_2282 + _GEN_1186; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1187 = {{3'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2284 = _T_2283 + _GEN_1187; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1188 = {{4'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2285 = _T_2284 + _GEN_1188; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1189 = {{5'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2286 = _T_2285 + _GEN_1189; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1190 = {{6'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2287 = _T_2286 + _GEN_1190; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2288 = 8'h2 == _T_2287; // @[Conditional.scala 37:30]
  wire  _T_2290 = 8'h3 == _T_2287; // @[Conditional.scala 37:30]
  wire  _GEN_225 = _T_2288 ? regs[112] : _T_2290; // @[Conditional.scala 40:58]
  wire [1:0] _T_2299 = regs[96] + regs[97]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1191 = {{1'd0}, regs[98]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2300 = _T_2299 + _GEN_1191; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1192 = {{2'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2301 = _T_2300 + _GEN_1192; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1193 = {{3'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2302 = _T_2301 + _GEN_1193; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1194 = {{4'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2303 = _T_2302 + _GEN_1194; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1195 = {{5'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2304 = _T_2303 + _GEN_1195; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1196 = {{6'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2305 = _T_2304 + _GEN_1196; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2306 = 8'h2 == _T_2305; // @[Conditional.scala 37:30]
  wire  _T_2308 = 8'h3 == _T_2305; // @[Conditional.scala 37:30]
  wire  _GEN_227 = _T_2306 ? regs[113] : _T_2308; // @[Conditional.scala 40:58]
  wire [1:0] _T_2317 = regs[97] + regs[98]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1197 = {{1'd0}, regs[99]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2318 = _T_2317 + _GEN_1197; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1198 = {{2'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2319 = _T_2318 + _GEN_1198; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1199 = {{3'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2320 = _T_2319 + _GEN_1199; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1200 = {{4'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2321 = _T_2320 + _GEN_1200; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1201 = {{5'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2322 = _T_2321 + _GEN_1201; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1202 = {{6'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2323 = _T_2322 + _GEN_1202; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2324 = 8'h2 == _T_2323; // @[Conditional.scala 37:30]
  wire  _T_2326 = 8'h3 == _T_2323; // @[Conditional.scala 37:30]
  wire  _GEN_229 = _T_2324 ? regs[114] : _T_2326; // @[Conditional.scala 40:58]
  wire [1:0] _T_2335 = regs[98] + regs[99]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1203 = {{1'd0}, regs[100]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2336 = _T_2335 + _GEN_1203; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1204 = {{2'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2337 = _T_2336 + _GEN_1204; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1205 = {{3'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2338 = _T_2337 + _GEN_1205; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1206 = {{4'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2339 = _T_2338 + _GEN_1206; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1207 = {{5'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2340 = _T_2339 + _GEN_1207; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1208 = {{6'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2341 = _T_2340 + _GEN_1208; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2342 = 8'h2 == _T_2341; // @[Conditional.scala 37:30]
  wire  _T_2344 = 8'h3 == _T_2341; // @[Conditional.scala 37:30]
  wire  _GEN_231 = _T_2342 ? regs[115] : _T_2344; // @[Conditional.scala 40:58]
  wire [1:0] _T_2353 = regs[99] + regs[100]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1209 = {{1'd0}, regs[101]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2354 = _T_2353 + _GEN_1209; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1210 = {{2'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2355 = _T_2354 + _GEN_1210; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1211 = {{3'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2356 = _T_2355 + _GEN_1211; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1212 = {{4'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2357 = _T_2356 + _GEN_1212; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1213 = {{5'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2358 = _T_2357 + _GEN_1213; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1214 = {{6'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2359 = _T_2358 + _GEN_1214; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2360 = 8'h2 == _T_2359; // @[Conditional.scala 37:30]
  wire  _T_2362 = 8'h3 == _T_2359; // @[Conditional.scala 37:30]
  wire  _GEN_233 = _T_2360 ? regs[116] : _T_2362; // @[Conditional.scala 40:58]
  wire [1:0] _T_2371 = regs[100] + regs[101]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1215 = {{1'd0}, regs[102]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2372 = _T_2371 + _GEN_1215; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1216 = {{2'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2373 = _T_2372 + _GEN_1216; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1217 = {{3'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2374 = _T_2373 + _GEN_1217; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1218 = {{4'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2375 = _T_2374 + _GEN_1218; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1219 = {{5'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2376 = _T_2375 + _GEN_1219; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1220 = {{6'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2377 = _T_2376 + _GEN_1220; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2378 = 8'h2 == _T_2377; // @[Conditional.scala 37:30]
  wire  _T_2380 = 8'h3 == _T_2377; // @[Conditional.scala 37:30]
  wire  _GEN_235 = _T_2378 ? regs[117] : _T_2380; // @[Conditional.scala 40:58]
  wire [1:0] _T_2389 = regs[101] + regs[102]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1221 = {{1'd0}, regs[103]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2390 = _T_2389 + _GEN_1221; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1222 = {{2'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2391 = _T_2390 + _GEN_1222; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1223 = {{3'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2392 = _T_2391 + _GEN_1223; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1224 = {{4'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2393 = _T_2392 + _GEN_1224; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1225 = {{5'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2394 = _T_2393 + _GEN_1225; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1226 = {{6'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2395 = _T_2394 + _GEN_1226; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2396 = 8'h2 == _T_2395; // @[Conditional.scala 37:30]
  wire  _T_2398 = 8'h3 == _T_2395; // @[Conditional.scala 37:30]
  wire  _GEN_237 = _T_2396 ? regs[118] : _T_2398; // @[Conditional.scala 40:58]
  wire [1:0] _T_2407 = regs[102] + regs[103]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1227 = {{1'd0}, regs[104]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2408 = _T_2407 + _GEN_1227; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1228 = {{2'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2409 = _T_2408 + _GEN_1228; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1229 = {{3'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2410 = _T_2409 + _GEN_1229; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1230 = {{4'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2411 = _T_2410 + _GEN_1230; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1231 = {{5'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2412 = _T_2411 + _GEN_1231; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1232 = {{6'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2413 = _T_2412 + _GEN_1232; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2414 = 8'h2 == _T_2413; // @[Conditional.scala 37:30]
  wire  _T_2416 = 8'h3 == _T_2413; // @[Conditional.scala 37:30]
  wire  _GEN_239 = _T_2414 ? regs[119] : _T_2416; // @[Conditional.scala 40:58]
  wire [1:0] _T_2425 = regs[103] + regs[104]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1233 = {{1'd0}, regs[105]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2426 = _T_2425 + _GEN_1233; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1234 = {{2'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2427 = _T_2426 + _GEN_1234; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1235 = {{3'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2428 = _T_2427 + _GEN_1235; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1236 = {{4'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2429 = _T_2428 + _GEN_1236; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1237 = {{5'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2430 = _T_2429 + _GEN_1237; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1238 = {{6'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2431 = _T_2430 + _GEN_1238; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2432 = 8'h2 == _T_2431; // @[Conditional.scala 37:30]
  wire  _T_2434 = 8'h3 == _T_2431; // @[Conditional.scala 37:30]
  wire  _GEN_241 = _T_2432 ? regs[120] : _T_2434; // @[Conditional.scala 40:58]
  wire [1:0] _T_2443 = regs[104] + regs[105]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1239 = {{1'd0}, regs[106]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2444 = _T_2443 + _GEN_1239; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1240 = {{2'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2445 = _T_2444 + _GEN_1240; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1241 = {{3'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2446 = _T_2445 + _GEN_1241; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1242 = {{4'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2447 = _T_2446 + _GEN_1242; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1243 = {{5'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2448 = _T_2447 + _GEN_1243; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1244 = {{6'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2449 = _T_2448 + _GEN_1244; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2450 = 8'h2 == _T_2449; // @[Conditional.scala 37:30]
  wire  _T_2452 = 8'h3 == _T_2449; // @[Conditional.scala 37:30]
  wire  _GEN_243 = _T_2450 ? regs[121] : _T_2452; // @[Conditional.scala 40:58]
  wire [1:0] _T_2461 = regs[105] + regs[106]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1245 = {{1'd0}, regs[107]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2462 = _T_2461 + _GEN_1245; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1246 = {{2'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2463 = _T_2462 + _GEN_1246; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1247 = {{3'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2464 = _T_2463 + _GEN_1247; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1248 = {{4'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2465 = _T_2464 + _GEN_1248; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1249 = {{5'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2466 = _T_2465 + _GEN_1249; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1250 = {{6'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2467 = _T_2466 + _GEN_1250; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2468 = 8'h2 == _T_2467; // @[Conditional.scala 37:30]
  wire  _T_2470 = 8'h3 == _T_2467; // @[Conditional.scala 37:30]
  wire  _GEN_245 = _T_2468 ? regs[122] : _T_2470; // @[Conditional.scala 40:58]
  wire [1:0] _T_2479 = regs[106] + regs[107]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1251 = {{1'd0}, regs[108]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2480 = _T_2479 + _GEN_1251; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1252 = {{2'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2481 = _T_2480 + _GEN_1252; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1253 = {{3'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2482 = _T_2481 + _GEN_1253; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1254 = {{4'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2483 = _T_2482 + _GEN_1254; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1255 = {{5'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2484 = _T_2483 + _GEN_1255; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1256 = {{6'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2485 = _T_2484 + _GEN_1256; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2486 = 8'h2 == _T_2485; // @[Conditional.scala 37:30]
  wire  _T_2488 = 8'h3 == _T_2485; // @[Conditional.scala 37:30]
  wire  _GEN_247 = _T_2486 ? regs[123] : _T_2488; // @[Conditional.scala 40:58]
  wire [1:0] _T_2497 = regs[107] + regs[108]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1257 = {{1'd0}, regs[109]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2498 = _T_2497 + _GEN_1257; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1258 = {{2'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2499 = _T_2498 + _GEN_1258; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1259 = {{3'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2500 = _T_2499 + _GEN_1259; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1260 = {{4'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2501 = _T_2500 + _GEN_1260; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1261 = {{5'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2502 = _T_2501 + _GEN_1261; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1262 = {{6'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2503 = _T_2502 + _GEN_1262; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2504 = 8'h2 == _T_2503; // @[Conditional.scala 37:30]
  wire  _T_2506 = 8'h3 == _T_2503; // @[Conditional.scala 37:30]
  wire  _GEN_249 = _T_2504 ? regs[124] : _T_2506; // @[Conditional.scala 40:58]
  wire [1:0] _T_2515 = regs[108] + regs[109]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1263 = {{1'd0}, regs[110]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2516 = _T_2515 + _GEN_1263; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1264 = {{2'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2517 = _T_2516 + _GEN_1264; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1265 = {{3'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2518 = _T_2517 + _GEN_1265; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1266 = {{4'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2519 = _T_2518 + _GEN_1266; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1267 = {{5'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2520 = _T_2519 + _GEN_1267; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1268 = {{6'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2521 = _T_2520 + _GEN_1268; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2522 = 8'h2 == _T_2521; // @[Conditional.scala 37:30]
  wire  _T_2524 = 8'h3 == _T_2521; // @[Conditional.scala 37:30]
  wire  _GEN_251 = _T_2522 ? regs[125] : _T_2524; // @[Conditional.scala 40:58]
  wire [1:0] _T_2533 = regs[109] + regs[110]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1269 = {{1'd0}, regs[111]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2534 = _T_2533 + _GEN_1269; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1270 = {{2'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2535 = _T_2534 + _GEN_1270; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1271 = {{3'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2536 = _T_2535 + _GEN_1271; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1272 = {{4'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2537 = _T_2536 + _GEN_1272; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1273 = {{5'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2538 = _T_2537 + _GEN_1273; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1274 = {{6'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2539 = _T_2538 + _GEN_1274; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2540 = 8'h2 == _T_2539; // @[Conditional.scala 37:30]
  wire  _T_2542 = 8'h3 == _T_2539; // @[Conditional.scala 37:30]
  wire  _GEN_253 = _T_2540 ? regs[126] : _T_2542; // @[Conditional.scala 40:58]
  wire [1:0] _T_2551 = regs[110] + regs[111]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1275 = {{1'd0}, regs[96]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2552 = _T_2551 + _GEN_1275; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1276 = {{2'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2553 = _T_2552 + _GEN_1276; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1277 = {{3'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2554 = _T_2553 + _GEN_1277; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1278 = {{4'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2555 = _T_2554 + _GEN_1278; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1279 = {{5'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2556 = _T_2555 + _GEN_1279; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1280 = {{6'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2557 = _T_2556 + _GEN_1280; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2558 = 8'h2 == _T_2557; // @[Conditional.scala 37:30]
  wire  _T_2560 = 8'h3 == _T_2557; // @[Conditional.scala 37:30]
  wire  _GEN_255 = _T_2558 ? regs[127] : _T_2560; // @[Conditional.scala 40:58]
  wire [1:0] _T_2569 = regs[127] + regs[112]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1281 = {{1'd0}, regs[113]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2570 = _T_2569 + _GEN_1281; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1282 = {{2'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2571 = _T_2570 + _GEN_1282; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1283 = {{3'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2572 = _T_2571 + _GEN_1283; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1284 = {{4'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2573 = _T_2572 + _GEN_1284; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1285 = {{5'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2574 = _T_2573 + _GEN_1285; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1286 = {{6'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2575 = _T_2574 + _GEN_1286; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2576 = 8'h2 == _T_2575; // @[Conditional.scala 37:30]
  wire  _T_2578 = 8'h3 == _T_2575; // @[Conditional.scala 37:30]
  wire  _GEN_257 = _T_2576 ? regs[128] : _T_2578; // @[Conditional.scala 40:58]
  wire [1:0] _T_2587 = regs[112] + regs[113]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1287 = {{1'd0}, regs[114]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2588 = _T_2587 + _GEN_1287; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1288 = {{2'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2589 = _T_2588 + _GEN_1288; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1289 = {{3'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2590 = _T_2589 + _GEN_1289; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1290 = {{4'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2591 = _T_2590 + _GEN_1290; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1291 = {{5'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2592 = _T_2591 + _GEN_1291; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1292 = {{6'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2593 = _T_2592 + _GEN_1292; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2594 = 8'h2 == _T_2593; // @[Conditional.scala 37:30]
  wire  _T_2596 = 8'h3 == _T_2593; // @[Conditional.scala 37:30]
  wire  _GEN_259 = _T_2594 ? regs[129] : _T_2596; // @[Conditional.scala 40:58]
  wire [1:0] _T_2605 = regs[113] + regs[114]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1293 = {{1'd0}, regs[115]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2606 = _T_2605 + _GEN_1293; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1294 = {{2'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2607 = _T_2606 + _GEN_1294; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1295 = {{3'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2608 = _T_2607 + _GEN_1295; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1296 = {{4'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2609 = _T_2608 + _GEN_1296; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1297 = {{5'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2610 = _T_2609 + _GEN_1297; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1298 = {{6'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2611 = _T_2610 + _GEN_1298; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2612 = 8'h2 == _T_2611; // @[Conditional.scala 37:30]
  wire  _T_2614 = 8'h3 == _T_2611; // @[Conditional.scala 37:30]
  wire  _GEN_261 = _T_2612 ? regs[130] : _T_2614; // @[Conditional.scala 40:58]
  wire [1:0] _T_2623 = regs[114] + regs[115]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1299 = {{1'd0}, regs[116]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2624 = _T_2623 + _GEN_1299; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1300 = {{2'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2625 = _T_2624 + _GEN_1300; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1301 = {{3'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2626 = _T_2625 + _GEN_1301; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1302 = {{4'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2627 = _T_2626 + _GEN_1302; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1303 = {{5'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2628 = _T_2627 + _GEN_1303; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1304 = {{6'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2629 = _T_2628 + _GEN_1304; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2630 = 8'h2 == _T_2629; // @[Conditional.scala 37:30]
  wire  _T_2632 = 8'h3 == _T_2629; // @[Conditional.scala 37:30]
  wire  _GEN_263 = _T_2630 ? regs[131] : _T_2632; // @[Conditional.scala 40:58]
  wire [1:0] _T_2641 = regs[115] + regs[116]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1305 = {{1'd0}, regs[117]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2642 = _T_2641 + _GEN_1305; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1306 = {{2'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2643 = _T_2642 + _GEN_1306; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1307 = {{3'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2644 = _T_2643 + _GEN_1307; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1308 = {{4'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2645 = _T_2644 + _GEN_1308; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1309 = {{5'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2646 = _T_2645 + _GEN_1309; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1310 = {{6'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2647 = _T_2646 + _GEN_1310; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2648 = 8'h2 == _T_2647; // @[Conditional.scala 37:30]
  wire  _T_2650 = 8'h3 == _T_2647; // @[Conditional.scala 37:30]
  wire  _GEN_265 = _T_2648 ? regs[132] : _T_2650; // @[Conditional.scala 40:58]
  wire [1:0] _T_2659 = regs[116] + regs[117]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1311 = {{1'd0}, regs[118]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2660 = _T_2659 + _GEN_1311; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1312 = {{2'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2661 = _T_2660 + _GEN_1312; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1313 = {{3'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2662 = _T_2661 + _GEN_1313; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1314 = {{4'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2663 = _T_2662 + _GEN_1314; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1315 = {{5'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2664 = _T_2663 + _GEN_1315; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1316 = {{6'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2665 = _T_2664 + _GEN_1316; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2666 = 8'h2 == _T_2665; // @[Conditional.scala 37:30]
  wire  _T_2668 = 8'h3 == _T_2665; // @[Conditional.scala 37:30]
  wire  _GEN_267 = _T_2666 ? regs[133] : _T_2668; // @[Conditional.scala 40:58]
  wire [1:0] _T_2677 = regs[117] + regs[118]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1317 = {{1'd0}, regs[119]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2678 = _T_2677 + _GEN_1317; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1318 = {{2'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2679 = _T_2678 + _GEN_1318; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1319 = {{3'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2680 = _T_2679 + _GEN_1319; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1320 = {{4'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2681 = _T_2680 + _GEN_1320; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1321 = {{5'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2682 = _T_2681 + _GEN_1321; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1322 = {{6'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2683 = _T_2682 + _GEN_1322; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2684 = 8'h2 == _T_2683; // @[Conditional.scala 37:30]
  wire  _T_2686 = 8'h3 == _T_2683; // @[Conditional.scala 37:30]
  wire  _GEN_269 = _T_2684 ? regs[134] : _T_2686; // @[Conditional.scala 40:58]
  wire [1:0] _T_2695 = regs[118] + regs[119]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1323 = {{1'd0}, regs[120]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2696 = _T_2695 + _GEN_1323; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1324 = {{2'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2697 = _T_2696 + _GEN_1324; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1325 = {{3'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2698 = _T_2697 + _GEN_1325; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1326 = {{4'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2699 = _T_2698 + _GEN_1326; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1327 = {{5'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2700 = _T_2699 + _GEN_1327; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1328 = {{6'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2701 = _T_2700 + _GEN_1328; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2702 = 8'h2 == _T_2701; // @[Conditional.scala 37:30]
  wire  _T_2704 = 8'h3 == _T_2701; // @[Conditional.scala 37:30]
  wire  _GEN_271 = _T_2702 ? regs[135] : _T_2704; // @[Conditional.scala 40:58]
  wire [1:0] _T_2713 = regs[119] + regs[120]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1329 = {{1'd0}, regs[121]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2714 = _T_2713 + _GEN_1329; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1330 = {{2'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2715 = _T_2714 + _GEN_1330; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1331 = {{3'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2716 = _T_2715 + _GEN_1331; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1332 = {{4'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2717 = _T_2716 + _GEN_1332; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1333 = {{5'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2718 = _T_2717 + _GEN_1333; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1334 = {{6'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2719 = _T_2718 + _GEN_1334; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2720 = 8'h2 == _T_2719; // @[Conditional.scala 37:30]
  wire  _T_2722 = 8'h3 == _T_2719; // @[Conditional.scala 37:30]
  wire  _GEN_273 = _T_2720 ? regs[136] : _T_2722; // @[Conditional.scala 40:58]
  wire [1:0] _T_2731 = regs[120] + regs[121]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1335 = {{1'd0}, regs[122]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2732 = _T_2731 + _GEN_1335; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1336 = {{2'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2733 = _T_2732 + _GEN_1336; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1337 = {{3'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2734 = _T_2733 + _GEN_1337; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1338 = {{4'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2735 = _T_2734 + _GEN_1338; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1339 = {{5'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2736 = _T_2735 + _GEN_1339; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1340 = {{6'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2737 = _T_2736 + _GEN_1340; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2738 = 8'h2 == _T_2737; // @[Conditional.scala 37:30]
  wire  _T_2740 = 8'h3 == _T_2737; // @[Conditional.scala 37:30]
  wire  _GEN_275 = _T_2738 ? regs[137] : _T_2740; // @[Conditional.scala 40:58]
  wire [1:0] _T_2749 = regs[121] + regs[122]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1341 = {{1'd0}, regs[123]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2750 = _T_2749 + _GEN_1341; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1342 = {{2'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2751 = _T_2750 + _GEN_1342; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1343 = {{3'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2752 = _T_2751 + _GEN_1343; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1344 = {{4'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2753 = _T_2752 + _GEN_1344; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1345 = {{5'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2754 = _T_2753 + _GEN_1345; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1346 = {{6'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2755 = _T_2754 + _GEN_1346; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2756 = 8'h2 == _T_2755; // @[Conditional.scala 37:30]
  wire  _T_2758 = 8'h3 == _T_2755; // @[Conditional.scala 37:30]
  wire  _GEN_277 = _T_2756 ? regs[138] : _T_2758; // @[Conditional.scala 40:58]
  wire [1:0] _T_2767 = regs[122] + regs[123]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1347 = {{1'd0}, regs[124]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2768 = _T_2767 + _GEN_1347; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1348 = {{2'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2769 = _T_2768 + _GEN_1348; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1349 = {{3'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2770 = _T_2769 + _GEN_1349; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1350 = {{4'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2771 = _T_2770 + _GEN_1350; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1351 = {{5'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2772 = _T_2771 + _GEN_1351; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1352 = {{6'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2773 = _T_2772 + _GEN_1352; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2774 = 8'h2 == _T_2773; // @[Conditional.scala 37:30]
  wire  _T_2776 = 8'h3 == _T_2773; // @[Conditional.scala 37:30]
  wire  _GEN_279 = _T_2774 ? regs[139] : _T_2776; // @[Conditional.scala 40:58]
  wire [1:0] _T_2785 = regs[123] + regs[124]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1353 = {{1'd0}, regs[125]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2786 = _T_2785 + _GEN_1353; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1354 = {{2'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2787 = _T_2786 + _GEN_1354; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1355 = {{3'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2788 = _T_2787 + _GEN_1355; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1356 = {{4'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2789 = _T_2788 + _GEN_1356; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1357 = {{5'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2790 = _T_2789 + _GEN_1357; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1358 = {{6'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2791 = _T_2790 + _GEN_1358; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2792 = 8'h2 == _T_2791; // @[Conditional.scala 37:30]
  wire  _T_2794 = 8'h3 == _T_2791; // @[Conditional.scala 37:30]
  wire  _GEN_281 = _T_2792 ? regs[140] : _T_2794; // @[Conditional.scala 40:58]
  wire [1:0] _T_2803 = regs[124] + regs[125]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1359 = {{1'd0}, regs[126]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2804 = _T_2803 + _GEN_1359; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1360 = {{2'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2805 = _T_2804 + _GEN_1360; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1361 = {{3'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2806 = _T_2805 + _GEN_1361; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1362 = {{4'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2807 = _T_2806 + _GEN_1362; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1363 = {{5'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2808 = _T_2807 + _GEN_1363; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1364 = {{6'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2809 = _T_2808 + _GEN_1364; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2810 = 8'h2 == _T_2809; // @[Conditional.scala 37:30]
  wire  _T_2812 = 8'h3 == _T_2809; // @[Conditional.scala 37:30]
  wire  _GEN_283 = _T_2810 ? regs[141] : _T_2812; // @[Conditional.scala 40:58]
  wire [1:0] _T_2821 = regs[125] + regs[126]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1365 = {{1'd0}, regs[127]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2822 = _T_2821 + _GEN_1365; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1366 = {{2'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2823 = _T_2822 + _GEN_1366; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1367 = {{3'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2824 = _T_2823 + _GEN_1367; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1368 = {{4'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2825 = _T_2824 + _GEN_1368; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1369 = {{5'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2826 = _T_2825 + _GEN_1369; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1370 = {{6'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2827 = _T_2826 + _GEN_1370; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2828 = 8'h2 == _T_2827; // @[Conditional.scala 37:30]
  wire  _T_2830 = 8'h3 == _T_2827; // @[Conditional.scala 37:30]
  wire  _GEN_285 = _T_2828 ? regs[142] : _T_2830; // @[Conditional.scala 40:58]
  wire [1:0] _T_2839 = regs[126] + regs[127]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1371 = {{1'd0}, regs[112]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2840 = _T_2839 + _GEN_1371; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1372 = {{2'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2841 = _T_2840 + _GEN_1372; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1373 = {{3'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2842 = _T_2841 + _GEN_1373; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1374 = {{4'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2843 = _T_2842 + _GEN_1374; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1375 = {{5'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2844 = _T_2843 + _GEN_1375; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1376 = {{6'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2845 = _T_2844 + _GEN_1376; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2846 = 8'h2 == _T_2845; // @[Conditional.scala 37:30]
  wire  _T_2848 = 8'h3 == _T_2845; // @[Conditional.scala 37:30]
  wire  _GEN_287 = _T_2846 ? regs[143] : _T_2848; // @[Conditional.scala 40:58]
  wire [1:0] _T_2857 = regs[143] + regs[128]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1377 = {{1'd0}, regs[129]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2858 = _T_2857 + _GEN_1377; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1378 = {{2'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2859 = _T_2858 + _GEN_1378; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1379 = {{3'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2860 = _T_2859 + _GEN_1379; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1380 = {{4'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2861 = _T_2860 + _GEN_1380; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1381 = {{5'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2862 = _T_2861 + _GEN_1381; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1382 = {{6'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2863 = _T_2862 + _GEN_1382; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2864 = 8'h2 == _T_2863; // @[Conditional.scala 37:30]
  wire  _T_2866 = 8'h3 == _T_2863; // @[Conditional.scala 37:30]
  wire  _GEN_289 = _T_2864 ? regs[144] : _T_2866; // @[Conditional.scala 40:58]
  wire [1:0] _T_2875 = regs[128] + regs[129]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1383 = {{1'd0}, regs[130]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2876 = _T_2875 + _GEN_1383; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1384 = {{2'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2877 = _T_2876 + _GEN_1384; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1385 = {{3'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2878 = _T_2877 + _GEN_1385; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1386 = {{4'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2879 = _T_2878 + _GEN_1386; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1387 = {{5'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2880 = _T_2879 + _GEN_1387; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1388 = {{6'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2881 = _T_2880 + _GEN_1388; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2882 = 8'h2 == _T_2881; // @[Conditional.scala 37:30]
  wire  _T_2884 = 8'h3 == _T_2881; // @[Conditional.scala 37:30]
  wire  _GEN_291 = _T_2882 ? regs[145] : _T_2884; // @[Conditional.scala 40:58]
  wire [1:0] _T_2893 = regs[129] + regs[130]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1389 = {{1'd0}, regs[131]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2894 = _T_2893 + _GEN_1389; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1390 = {{2'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2895 = _T_2894 + _GEN_1390; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1391 = {{3'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2896 = _T_2895 + _GEN_1391; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1392 = {{4'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2897 = _T_2896 + _GEN_1392; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1393 = {{5'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2898 = _T_2897 + _GEN_1393; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1394 = {{6'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2899 = _T_2898 + _GEN_1394; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2900 = 8'h2 == _T_2899; // @[Conditional.scala 37:30]
  wire  _T_2902 = 8'h3 == _T_2899; // @[Conditional.scala 37:30]
  wire  _GEN_293 = _T_2900 ? regs[146] : _T_2902; // @[Conditional.scala 40:58]
  wire [1:0] _T_2911 = regs[130] + regs[131]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1395 = {{1'd0}, regs[132]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2912 = _T_2911 + _GEN_1395; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1396 = {{2'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2913 = _T_2912 + _GEN_1396; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1397 = {{3'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2914 = _T_2913 + _GEN_1397; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1398 = {{4'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2915 = _T_2914 + _GEN_1398; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1399 = {{5'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2916 = _T_2915 + _GEN_1399; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1400 = {{6'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2917 = _T_2916 + _GEN_1400; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2918 = 8'h2 == _T_2917; // @[Conditional.scala 37:30]
  wire  _T_2920 = 8'h3 == _T_2917; // @[Conditional.scala 37:30]
  wire  _GEN_295 = _T_2918 ? regs[147] : _T_2920; // @[Conditional.scala 40:58]
  wire [1:0] _T_2929 = regs[131] + regs[132]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1401 = {{1'd0}, regs[133]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2930 = _T_2929 + _GEN_1401; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1402 = {{2'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2931 = _T_2930 + _GEN_1402; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1403 = {{3'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2932 = _T_2931 + _GEN_1403; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1404 = {{4'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2933 = _T_2932 + _GEN_1404; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1405 = {{5'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2934 = _T_2933 + _GEN_1405; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1406 = {{6'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2935 = _T_2934 + _GEN_1406; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2936 = 8'h2 == _T_2935; // @[Conditional.scala 37:30]
  wire  _T_2938 = 8'h3 == _T_2935; // @[Conditional.scala 37:30]
  wire  _GEN_297 = _T_2936 ? regs[148] : _T_2938; // @[Conditional.scala 40:58]
  wire [1:0] _T_2947 = regs[132] + regs[133]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1407 = {{1'd0}, regs[134]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2948 = _T_2947 + _GEN_1407; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1408 = {{2'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2949 = _T_2948 + _GEN_1408; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1409 = {{3'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2950 = _T_2949 + _GEN_1409; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1410 = {{4'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2951 = _T_2950 + _GEN_1410; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1411 = {{5'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2952 = _T_2951 + _GEN_1411; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1412 = {{6'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2953 = _T_2952 + _GEN_1412; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2954 = 8'h2 == _T_2953; // @[Conditional.scala 37:30]
  wire  _T_2956 = 8'h3 == _T_2953; // @[Conditional.scala 37:30]
  wire  _GEN_299 = _T_2954 ? regs[149] : _T_2956; // @[Conditional.scala 40:58]
  wire [1:0] _T_2965 = regs[133] + regs[134]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1413 = {{1'd0}, regs[135]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2966 = _T_2965 + _GEN_1413; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1414 = {{2'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2967 = _T_2966 + _GEN_1414; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1415 = {{3'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2968 = _T_2967 + _GEN_1415; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1416 = {{4'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2969 = _T_2968 + _GEN_1416; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1417 = {{5'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2970 = _T_2969 + _GEN_1417; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1418 = {{6'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2971 = _T_2970 + _GEN_1418; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2972 = 8'h2 == _T_2971; // @[Conditional.scala 37:30]
  wire  _T_2974 = 8'h3 == _T_2971; // @[Conditional.scala 37:30]
  wire  _GEN_301 = _T_2972 ? regs[150] : _T_2974; // @[Conditional.scala 40:58]
  wire [1:0] _T_2983 = regs[134] + regs[135]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1419 = {{1'd0}, regs[136]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_2984 = _T_2983 + _GEN_1419; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1420 = {{2'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_2985 = _T_2984 + _GEN_1420; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1421 = {{3'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_2986 = _T_2985 + _GEN_1421; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1422 = {{4'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_2987 = _T_2986 + _GEN_1422; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1423 = {{5'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_2988 = _T_2987 + _GEN_1423; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1424 = {{6'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_2989 = _T_2988 + _GEN_1424; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_2990 = 8'h2 == _T_2989; // @[Conditional.scala 37:30]
  wire  _T_2992 = 8'h3 == _T_2989; // @[Conditional.scala 37:30]
  wire  _GEN_303 = _T_2990 ? regs[151] : _T_2992; // @[Conditional.scala 40:58]
  wire [1:0] _T_3001 = regs[135] + regs[136]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1425 = {{1'd0}, regs[137]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3002 = _T_3001 + _GEN_1425; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1426 = {{2'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3003 = _T_3002 + _GEN_1426; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1427 = {{3'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3004 = _T_3003 + _GEN_1427; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1428 = {{4'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3005 = _T_3004 + _GEN_1428; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1429 = {{5'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3006 = _T_3005 + _GEN_1429; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1430 = {{6'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3007 = _T_3006 + _GEN_1430; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3008 = 8'h2 == _T_3007; // @[Conditional.scala 37:30]
  wire  _T_3010 = 8'h3 == _T_3007; // @[Conditional.scala 37:30]
  wire  _GEN_305 = _T_3008 ? regs[152] : _T_3010; // @[Conditional.scala 40:58]
  wire [1:0] _T_3019 = regs[136] + regs[137]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1431 = {{1'd0}, regs[138]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3020 = _T_3019 + _GEN_1431; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1432 = {{2'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3021 = _T_3020 + _GEN_1432; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1433 = {{3'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3022 = _T_3021 + _GEN_1433; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1434 = {{4'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3023 = _T_3022 + _GEN_1434; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1435 = {{5'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3024 = _T_3023 + _GEN_1435; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1436 = {{6'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3025 = _T_3024 + _GEN_1436; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3026 = 8'h2 == _T_3025; // @[Conditional.scala 37:30]
  wire  _T_3028 = 8'h3 == _T_3025; // @[Conditional.scala 37:30]
  wire  _GEN_307 = _T_3026 ? regs[153] : _T_3028; // @[Conditional.scala 40:58]
  wire [1:0] _T_3037 = regs[137] + regs[138]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1437 = {{1'd0}, regs[139]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3038 = _T_3037 + _GEN_1437; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1438 = {{2'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3039 = _T_3038 + _GEN_1438; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1439 = {{3'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3040 = _T_3039 + _GEN_1439; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1440 = {{4'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3041 = _T_3040 + _GEN_1440; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1441 = {{5'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3042 = _T_3041 + _GEN_1441; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1442 = {{6'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3043 = _T_3042 + _GEN_1442; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3044 = 8'h2 == _T_3043; // @[Conditional.scala 37:30]
  wire  _T_3046 = 8'h3 == _T_3043; // @[Conditional.scala 37:30]
  wire  _GEN_309 = _T_3044 ? regs[154] : _T_3046; // @[Conditional.scala 40:58]
  wire [1:0] _T_3055 = regs[138] + regs[139]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1443 = {{1'd0}, regs[140]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3056 = _T_3055 + _GEN_1443; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1444 = {{2'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3057 = _T_3056 + _GEN_1444; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1445 = {{3'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3058 = _T_3057 + _GEN_1445; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1446 = {{4'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3059 = _T_3058 + _GEN_1446; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1447 = {{5'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3060 = _T_3059 + _GEN_1447; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1448 = {{6'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3061 = _T_3060 + _GEN_1448; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3062 = 8'h2 == _T_3061; // @[Conditional.scala 37:30]
  wire  _T_3064 = 8'h3 == _T_3061; // @[Conditional.scala 37:30]
  wire  _GEN_311 = _T_3062 ? regs[155] : _T_3064; // @[Conditional.scala 40:58]
  wire [1:0] _T_3073 = regs[139] + regs[140]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1449 = {{1'd0}, regs[141]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3074 = _T_3073 + _GEN_1449; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1450 = {{2'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3075 = _T_3074 + _GEN_1450; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1451 = {{3'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3076 = _T_3075 + _GEN_1451; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1452 = {{4'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3077 = _T_3076 + _GEN_1452; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1453 = {{5'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3078 = _T_3077 + _GEN_1453; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1454 = {{6'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3079 = _T_3078 + _GEN_1454; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3080 = 8'h2 == _T_3079; // @[Conditional.scala 37:30]
  wire  _T_3082 = 8'h3 == _T_3079; // @[Conditional.scala 37:30]
  wire  _GEN_313 = _T_3080 ? regs[156] : _T_3082; // @[Conditional.scala 40:58]
  wire [1:0] _T_3091 = regs[140] + regs[141]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1455 = {{1'd0}, regs[142]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3092 = _T_3091 + _GEN_1455; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1456 = {{2'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3093 = _T_3092 + _GEN_1456; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1457 = {{3'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3094 = _T_3093 + _GEN_1457; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1458 = {{4'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3095 = _T_3094 + _GEN_1458; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1459 = {{5'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3096 = _T_3095 + _GEN_1459; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1460 = {{6'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3097 = _T_3096 + _GEN_1460; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3098 = 8'h2 == _T_3097; // @[Conditional.scala 37:30]
  wire  _T_3100 = 8'h3 == _T_3097; // @[Conditional.scala 37:30]
  wire  _GEN_315 = _T_3098 ? regs[157] : _T_3100; // @[Conditional.scala 40:58]
  wire [1:0] _T_3109 = regs[141] + regs[142]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1461 = {{1'd0}, regs[143]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3110 = _T_3109 + _GEN_1461; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1462 = {{2'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3111 = _T_3110 + _GEN_1462; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1463 = {{3'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3112 = _T_3111 + _GEN_1463; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1464 = {{4'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3113 = _T_3112 + _GEN_1464; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1465 = {{5'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3114 = _T_3113 + _GEN_1465; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1466 = {{6'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3115 = _T_3114 + _GEN_1466; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3116 = 8'h2 == _T_3115; // @[Conditional.scala 37:30]
  wire  _T_3118 = 8'h3 == _T_3115; // @[Conditional.scala 37:30]
  wire  _GEN_317 = _T_3116 ? regs[158] : _T_3118; // @[Conditional.scala 40:58]
  wire [1:0] _T_3127 = regs[142] + regs[143]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1467 = {{1'd0}, regs[128]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3128 = _T_3127 + _GEN_1467; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1468 = {{2'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3129 = _T_3128 + _GEN_1468; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1469 = {{3'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3130 = _T_3129 + _GEN_1469; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1470 = {{4'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3131 = _T_3130 + _GEN_1470; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1471 = {{5'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3132 = _T_3131 + _GEN_1471; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1472 = {{6'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3133 = _T_3132 + _GEN_1472; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3134 = 8'h2 == _T_3133; // @[Conditional.scala 37:30]
  wire  _T_3136 = 8'h3 == _T_3133; // @[Conditional.scala 37:30]
  wire  _GEN_319 = _T_3134 ? regs[159] : _T_3136; // @[Conditional.scala 40:58]
  wire [1:0] _T_3145 = regs[159] + regs[144]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1473 = {{1'd0}, regs[145]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3146 = _T_3145 + _GEN_1473; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1474 = {{2'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3147 = _T_3146 + _GEN_1474; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1475 = {{3'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3148 = _T_3147 + _GEN_1475; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1476 = {{4'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3149 = _T_3148 + _GEN_1476; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1477 = {{5'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3150 = _T_3149 + _GEN_1477; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1478 = {{6'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3151 = _T_3150 + _GEN_1478; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3152 = 8'h2 == _T_3151; // @[Conditional.scala 37:30]
  wire  _T_3154 = 8'h3 == _T_3151; // @[Conditional.scala 37:30]
  wire  _GEN_321 = _T_3152 ? regs[160] : _T_3154; // @[Conditional.scala 40:58]
  wire [1:0] _T_3163 = regs[144] + regs[145]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1479 = {{1'd0}, regs[146]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3164 = _T_3163 + _GEN_1479; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1480 = {{2'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3165 = _T_3164 + _GEN_1480; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1481 = {{3'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3166 = _T_3165 + _GEN_1481; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1482 = {{4'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3167 = _T_3166 + _GEN_1482; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1483 = {{5'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3168 = _T_3167 + _GEN_1483; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1484 = {{6'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3169 = _T_3168 + _GEN_1484; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3170 = 8'h2 == _T_3169; // @[Conditional.scala 37:30]
  wire  _T_3172 = 8'h3 == _T_3169; // @[Conditional.scala 37:30]
  wire  _GEN_323 = _T_3170 ? regs[161] : _T_3172; // @[Conditional.scala 40:58]
  wire [1:0] _T_3181 = regs[145] + regs[146]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1485 = {{1'd0}, regs[147]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3182 = _T_3181 + _GEN_1485; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1486 = {{2'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3183 = _T_3182 + _GEN_1486; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1487 = {{3'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3184 = _T_3183 + _GEN_1487; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1488 = {{4'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3185 = _T_3184 + _GEN_1488; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1489 = {{5'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3186 = _T_3185 + _GEN_1489; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1490 = {{6'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3187 = _T_3186 + _GEN_1490; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3188 = 8'h2 == _T_3187; // @[Conditional.scala 37:30]
  wire  _T_3190 = 8'h3 == _T_3187; // @[Conditional.scala 37:30]
  wire  _GEN_325 = _T_3188 ? regs[162] : _T_3190; // @[Conditional.scala 40:58]
  wire [1:0] _T_3199 = regs[146] + regs[147]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1491 = {{1'd0}, regs[148]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3200 = _T_3199 + _GEN_1491; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1492 = {{2'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3201 = _T_3200 + _GEN_1492; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1493 = {{3'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3202 = _T_3201 + _GEN_1493; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1494 = {{4'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3203 = _T_3202 + _GEN_1494; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1495 = {{5'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3204 = _T_3203 + _GEN_1495; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1496 = {{6'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3205 = _T_3204 + _GEN_1496; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3206 = 8'h2 == _T_3205; // @[Conditional.scala 37:30]
  wire  _T_3208 = 8'h3 == _T_3205; // @[Conditional.scala 37:30]
  wire  _GEN_327 = _T_3206 ? regs[163] : _T_3208; // @[Conditional.scala 40:58]
  wire [1:0] _T_3217 = regs[147] + regs[148]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1497 = {{1'd0}, regs[149]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3218 = _T_3217 + _GEN_1497; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1498 = {{2'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3219 = _T_3218 + _GEN_1498; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1499 = {{3'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3220 = _T_3219 + _GEN_1499; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1500 = {{4'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3221 = _T_3220 + _GEN_1500; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1501 = {{5'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3222 = _T_3221 + _GEN_1501; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1502 = {{6'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3223 = _T_3222 + _GEN_1502; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3224 = 8'h2 == _T_3223; // @[Conditional.scala 37:30]
  wire  _T_3226 = 8'h3 == _T_3223; // @[Conditional.scala 37:30]
  wire  _GEN_329 = _T_3224 ? regs[164] : _T_3226; // @[Conditional.scala 40:58]
  wire [1:0] _T_3235 = regs[148] + regs[149]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1503 = {{1'd0}, regs[150]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3236 = _T_3235 + _GEN_1503; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1504 = {{2'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3237 = _T_3236 + _GEN_1504; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1505 = {{3'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3238 = _T_3237 + _GEN_1505; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1506 = {{4'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3239 = _T_3238 + _GEN_1506; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1507 = {{5'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3240 = _T_3239 + _GEN_1507; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1508 = {{6'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3241 = _T_3240 + _GEN_1508; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3242 = 8'h2 == _T_3241; // @[Conditional.scala 37:30]
  wire  _T_3244 = 8'h3 == _T_3241; // @[Conditional.scala 37:30]
  wire  _GEN_331 = _T_3242 ? regs[165] : _T_3244; // @[Conditional.scala 40:58]
  wire [1:0] _T_3253 = regs[149] + regs[150]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1509 = {{1'd0}, regs[151]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3254 = _T_3253 + _GEN_1509; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1510 = {{2'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3255 = _T_3254 + _GEN_1510; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1511 = {{3'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3256 = _T_3255 + _GEN_1511; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1512 = {{4'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3257 = _T_3256 + _GEN_1512; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1513 = {{5'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3258 = _T_3257 + _GEN_1513; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1514 = {{6'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3259 = _T_3258 + _GEN_1514; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3260 = 8'h2 == _T_3259; // @[Conditional.scala 37:30]
  wire  _T_3262 = 8'h3 == _T_3259; // @[Conditional.scala 37:30]
  wire  _GEN_333 = _T_3260 ? regs[166] : _T_3262; // @[Conditional.scala 40:58]
  wire [1:0] _T_3271 = regs[150] + regs[151]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1515 = {{1'd0}, regs[152]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3272 = _T_3271 + _GEN_1515; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1516 = {{2'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3273 = _T_3272 + _GEN_1516; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1517 = {{3'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3274 = _T_3273 + _GEN_1517; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1518 = {{4'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3275 = _T_3274 + _GEN_1518; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1519 = {{5'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3276 = _T_3275 + _GEN_1519; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1520 = {{6'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3277 = _T_3276 + _GEN_1520; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3278 = 8'h2 == _T_3277; // @[Conditional.scala 37:30]
  wire  _T_3280 = 8'h3 == _T_3277; // @[Conditional.scala 37:30]
  wire  _GEN_335 = _T_3278 ? regs[167] : _T_3280; // @[Conditional.scala 40:58]
  wire [1:0] _T_3289 = regs[151] + regs[152]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1521 = {{1'd0}, regs[153]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3290 = _T_3289 + _GEN_1521; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1522 = {{2'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3291 = _T_3290 + _GEN_1522; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1523 = {{3'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3292 = _T_3291 + _GEN_1523; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1524 = {{4'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3293 = _T_3292 + _GEN_1524; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1525 = {{5'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3294 = _T_3293 + _GEN_1525; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1526 = {{6'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3295 = _T_3294 + _GEN_1526; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3296 = 8'h2 == _T_3295; // @[Conditional.scala 37:30]
  wire  _T_3298 = 8'h3 == _T_3295; // @[Conditional.scala 37:30]
  wire  _GEN_337 = _T_3296 ? regs[168] : _T_3298; // @[Conditional.scala 40:58]
  wire [1:0] _T_3307 = regs[152] + regs[153]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1527 = {{1'd0}, regs[154]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3308 = _T_3307 + _GEN_1527; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1528 = {{2'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3309 = _T_3308 + _GEN_1528; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1529 = {{3'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3310 = _T_3309 + _GEN_1529; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1530 = {{4'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3311 = _T_3310 + _GEN_1530; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1531 = {{5'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3312 = _T_3311 + _GEN_1531; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1532 = {{6'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3313 = _T_3312 + _GEN_1532; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3314 = 8'h2 == _T_3313; // @[Conditional.scala 37:30]
  wire  _T_3316 = 8'h3 == _T_3313; // @[Conditional.scala 37:30]
  wire  _GEN_339 = _T_3314 ? regs[169] : _T_3316; // @[Conditional.scala 40:58]
  wire [1:0] _T_3325 = regs[153] + regs[154]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1533 = {{1'd0}, regs[155]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3326 = _T_3325 + _GEN_1533; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1534 = {{2'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3327 = _T_3326 + _GEN_1534; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1535 = {{3'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3328 = _T_3327 + _GEN_1535; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1536 = {{4'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3329 = _T_3328 + _GEN_1536; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1537 = {{5'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3330 = _T_3329 + _GEN_1537; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1538 = {{6'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3331 = _T_3330 + _GEN_1538; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3332 = 8'h2 == _T_3331; // @[Conditional.scala 37:30]
  wire  _T_3334 = 8'h3 == _T_3331; // @[Conditional.scala 37:30]
  wire  _GEN_341 = _T_3332 ? regs[170] : _T_3334; // @[Conditional.scala 40:58]
  wire [1:0] _T_3343 = regs[154] + regs[155]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1539 = {{1'd0}, regs[156]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3344 = _T_3343 + _GEN_1539; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1540 = {{2'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3345 = _T_3344 + _GEN_1540; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1541 = {{3'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3346 = _T_3345 + _GEN_1541; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1542 = {{4'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3347 = _T_3346 + _GEN_1542; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1543 = {{5'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3348 = _T_3347 + _GEN_1543; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1544 = {{6'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3349 = _T_3348 + _GEN_1544; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3350 = 8'h2 == _T_3349; // @[Conditional.scala 37:30]
  wire  _T_3352 = 8'h3 == _T_3349; // @[Conditional.scala 37:30]
  wire  _GEN_343 = _T_3350 ? regs[171] : _T_3352; // @[Conditional.scala 40:58]
  wire [1:0] _T_3361 = regs[155] + regs[156]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1545 = {{1'd0}, regs[157]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3362 = _T_3361 + _GEN_1545; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1546 = {{2'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3363 = _T_3362 + _GEN_1546; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1547 = {{3'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3364 = _T_3363 + _GEN_1547; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1548 = {{4'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3365 = _T_3364 + _GEN_1548; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1549 = {{5'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3366 = _T_3365 + _GEN_1549; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1550 = {{6'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3367 = _T_3366 + _GEN_1550; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3368 = 8'h2 == _T_3367; // @[Conditional.scala 37:30]
  wire  _T_3370 = 8'h3 == _T_3367; // @[Conditional.scala 37:30]
  wire  _GEN_345 = _T_3368 ? regs[172] : _T_3370; // @[Conditional.scala 40:58]
  wire [1:0] _T_3379 = regs[156] + regs[157]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1551 = {{1'd0}, regs[158]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3380 = _T_3379 + _GEN_1551; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1552 = {{2'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3381 = _T_3380 + _GEN_1552; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1553 = {{3'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3382 = _T_3381 + _GEN_1553; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1554 = {{4'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3383 = _T_3382 + _GEN_1554; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1555 = {{5'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3384 = _T_3383 + _GEN_1555; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1556 = {{6'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3385 = _T_3384 + _GEN_1556; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3386 = 8'h2 == _T_3385; // @[Conditional.scala 37:30]
  wire  _T_3388 = 8'h3 == _T_3385; // @[Conditional.scala 37:30]
  wire  _GEN_347 = _T_3386 ? regs[173] : _T_3388; // @[Conditional.scala 40:58]
  wire [1:0] _T_3397 = regs[157] + regs[158]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1557 = {{1'd0}, regs[159]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3398 = _T_3397 + _GEN_1557; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1558 = {{2'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3399 = _T_3398 + _GEN_1558; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1559 = {{3'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3400 = _T_3399 + _GEN_1559; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1560 = {{4'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3401 = _T_3400 + _GEN_1560; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1561 = {{5'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3402 = _T_3401 + _GEN_1561; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1562 = {{6'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3403 = _T_3402 + _GEN_1562; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3404 = 8'h2 == _T_3403; // @[Conditional.scala 37:30]
  wire  _T_3406 = 8'h3 == _T_3403; // @[Conditional.scala 37:30]
  wire  _GEN_349 = _T_3404 ? regs[174] : _T_3406; // @[Conditional.scala 40:58]
  wire [1:0] _T_3415 = regs[158] + regs[159]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1563 = {{1'd0}, regs[144]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3416 = _T_3415 + _GEN_1563; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1564 = {{2'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3417 = _T_3416 + _GEN_1564; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1565 = {{3'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3418 = _T_3417 + _GEN_1565; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1566 = {{4'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3419 = _T_3418 + _GEN_1566; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1567 = {{5'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3420 = _T_3419 + _GEN_1567; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1568 = {{6'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3421 = _T_3420 + _GEN_1568; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3422 = 8'h2 == _T_3421; // @[Conditional.scala 37:30]
  wire  _T_3424 = 8'h3 == _T_3421; // @[Conditional.scala 37:30]
  wire  _GEN_351 = _T_3422 ? regs[175] : _T_3424; // @[Conditional.scala 40:58]
  wire [1:0] _T_3433 = regs[175] + regs[160]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1569 = {{1'd0}, regs[161]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3434 = _T_3433 + _GEN_1569; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1570 = {{2'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3435 = _T_3434 + _GEN_1570; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1571 = {{3'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3436 = _T_3435 + _GEN_1571; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1572 = {{4'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3437 = _T_3436 + _GEN_1572; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1573 = {{5'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3438 = _T_3437 + _GEN_1573; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1574 = {{6'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3439 = _T_3438 + _GEN_1574; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3440 = 8'h2 == _T_3439; // @[Conditional.scala 37:30]
  wire  _T_3442 = 8'h3 == _T_3439; // @[Conditional.scala 37:30]
  wire  _GEN_353 = _T_3440 ? regs[176] : _T_3442; // @[Conditional.scala 40:58]
  wire [1:0] _T_3451 = regs[160] + regs[161]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1575 = {{1'd0}, regs[162]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3452 = _T_3451 + _GEN_1575; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1576 = {{2'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3453 = _T_3452 + _GEN_1576; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1577 = {{3'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3454 = _T_3453 + _GEN_1577; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1578 = {{4'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3455 = _T_3454 + _GEN_1578; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1579 = {{5'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3456 = _T_3455 + _GEN_1579; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1580 = {{6'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3457 = _T_3456 + _GEN_1580; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3458 = 8'h2 == _T_3457; // @[Conditional.scala 37:30]
  wire  _T_3460 = 8'h3 == _T_3457; // @[Conditional.scala 37:30]
  wire  _GEN_355 = _T_3458 ? regs[177] : _T_3460; // @[Conditional.scala 40:58]
  wire [1:0] _T_3469 = regs[161] + regs[162]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1581 = {{1'd0}, regs[163]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3470 = _T_3469 + _GEN_1581; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1582 = {{2'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3471 = _T_3470 + _GEN_1582; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1583 = {{3'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3472 = _T_3471 + _GEN_1583; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1584 = {{4'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3473 = _T_3472 + _GEN_1584; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1585 = {{5'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3474 = _T_3473 + _GEN_1585; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1586 = {{6'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3475 = _T_3474 + _GEN_1586; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3476 = 8'h2 == _T_3475; // @[Conditional.scala 37:30]
  wire  _T_3478 = 8'h3 == _T_3475; // @[Conditional.scala 37:30]
  wire  _GEN_357 = _T_3476 ? regs[178] : _T_3478; // @[Conditional.scala 40:58]
  wire [1:0] _T_3487 = regs[162] + regs[163]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1587 = {{1'd0}, regs[164]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3488 = _T_3487 + _GEN_1587; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1588 = {{2'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3489 = _T_3488 + _GEN_1588; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1589 = {{3'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3490 = _T_3489 + _GEN_1589; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1590 = {{4'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3491 = _T_3490 + _GEN_1590; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1591 = {{5'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3492 = _T_3491 + _GEN_1591; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1592 = {{6'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3493 = _T_3492 + _GEN_1592; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3494 = 8'h2 == _T_3493; // @[Conditional.scala 37:30]
  wire  _T_3496 = 8'h3 == _T_3493; // @[Conditional.scala 37:30]
  wire  _GEN_359 = _T_3494 ? regs[179] : _T_3496; // @[Conditional.scala 40:58]
  wire [1:0] _T_3505 = regs[163] + regs[164]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1593 = {{1'd0}, regs[165]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3506 = _T_3505 + _GEN_1593; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1594 = {{2'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3507 = _T_3506 + _GEN_1594; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1595 = {{3'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3508 = _T_3507 + _GEN_1595; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1596 = {{4'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3509 = _T_3508 + _GEN_1596; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1597 = {{5'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3510 = _T_3509 + _GEN_1597; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1598 = {{6'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3511 = _T_3510 + _GEN_1598; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3512 = 8'h2 == _T_3511; // @[Conditional.scala 37:30]
  wire  _T_3514 = 8'h3 == _T_3511; // @[Conditional.scala 37:30]
  wire  _GEN_361 = _T_3512 ? regs[180] : _T_3514; // @[Conditional.scala 40:58]
  wire [1:0] _T_3523 = regs[164] + regs[165]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1599 = {{1'd0}, regs[166]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3524 = _T_3523 + _GEN_1599; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1600 = {{2'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3525 = _T_3524 + _GEN_1600; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1601 = {{3'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3526 = _T_3525 + _GEN_1601; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1602 = {{4'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3527 = _T_3526 + _GEN_1602; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1603 = {{5'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3528 = _T_3527 + _GEN_1603; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1604 = {{6'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3529 = _T_3528 + _GEN_1604; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3530 = 8'h2 == _T_3529; // @[Conditional.scala 37:30]
  wire  _T_3532 = 8'h3 == _T_3529; // @[Conditional.scala 37:30]
  wire  _GEN_363 = _T_3530 ? regs[181] : _T_3532; // @[Conditional.scala 40:58]
  wire [1:0] _T_3541 = regs[165] + regs[166]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1605 = {{1'd0}, regs[167]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3542 = _T_3541 + _GEN_1605; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1606 = {{2'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3543 = _T_3542 + _GEN_1606; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1607 = {{3'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3544 = _T_3543 + _GEN_1607; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1608 = {{4'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3545 = _T_3544 + _GEN_1608; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1609 = {{5'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3546 = _T_3545 + _GEN_1609; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1610 = {{6'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3547 = _T_3546 + _GEN_1610; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3548 = 8'h2 == _T_3547; // @[Conditional.scala 37:30]
  wire  _T_3550 = 8'h3 == _T_3547; // @[Conditional.scala 37:30]
  wire  _GEN_365 = _T_3548 ? regs[182] : _T_3550; // @[Conditional.scala 40:58]
  wire [1:0] _T_3559 = regs[166] + regs[167]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1611 = {{1'd0}, regs[168]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3560 = _T_3559 + _GEN_1611; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1612 = {{2'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3561 = _T_3560 + _GEN_1612; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1613 = {{3'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3562 = _T_3561 + _GEN_1613; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1614 = {{4'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3563 = _T_3562 + _GEN_1614; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1615 = {{5'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3564 = _T_3563 + _GEN_1615; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1616 = {{6'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3565 = _T_3564 + _GEN_1616; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3566 = 8'h2 == _T_3565; // @[Conditional.scala 37:30]
  wire  _T_3568 = 8'h3 == _T_3565; // @[Conditional.scala 37:30]
  wire  _GEN_367 = _T_3566 ? regs[183] : _T_3568; // @[Conditional.scala 40:58]
  wire [1:0] _T_3577 = regs[167] + regs[168]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1617 = {{1'd0}, regs[169]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3578 = _T_3577 + _GEN_1617; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1618 = {{2'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3579 = _T_3578 + _GEN_1618; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1619 = {{3'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3580 = _T_3579 + _GEN_1619; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1620 = {{4'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3581 = _T_3580 + _GEN_1620; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1621 = {{5'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3582 = _T_3581 + _GEN_1621; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1622 = {{6'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3583 = _T_3582 + _GEN_1622; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3584 = 8'h2 == _T_3583; // @[Conditional.scala 37:30]
  wire  _T_3586 = 8'h3 == _T_3583; // @[Conditional.scala 37:30]
  wire  _GEN_369 = _T_3584 ? regs[184] : _T_3586; // @[Conditional.scala 40:58]
  wire [1:0] _T_3595 = regs[168] + regs[169]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1623 = {{1'd0}, regs[170]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3596 = _T_3595 + _GEN_1623; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1624 = {{2'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3597 = _T_3596 + _GEN_1624; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1625 = {{3'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3598 = _T_3597 + _GEN_1625; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1626 = {{4'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3599 = _T_3598 + _GEN_1626; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1627 = {{5'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3600 = _T_3599 + _GEN_1627; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1628 = {{6'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3601 = _T_3600 + _GEN_1628; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3602 = 8'h2 == _T_3601; // @[Conditional.scala 37:30]
  wire  _T_3604 = 8'h3 == _T_3601; // @[Conditional.scala 37:30]
  wire  _GEN_371 = _T_3602 ? regs[185] : _T_3604; // @[Conditional.scala 40:58]
  wire [1:0] _T_3613 = regs[169] + regs[170]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1629 = {{1'd0}, regs[171]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3614 = _T_3613 + _GEN_1629; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1630 = {{2'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3615 = _T_3614 + _GEN_1630; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1631 = {{3'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3616 = _T_3615 + _GEN_1631; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1632 = {{4'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3617 = _T_3616 + _GEN_1632; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1633 = {{5'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3618 = _T_3617 + _GEN_1633; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1634 = {{6'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3619 = _T_3618 + _GEN_1634; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3620 = 8'h2 == _T_3619; // @[Conditional.scala 37:30]
  wire  _T_3622 = 8'h3 == _T_3619; // @[Conditional.scala 37:30]
  wire  _GEN_373 = _T_3620 ? regs[186] : _T_3622; // @[Conditional.scala 40:58]
  wire [1:0] _T_3631 = regs[170] + regs[171]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1635 = {{1'd0}, regs[172]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3632 = _T_3631 + _GEN_1635; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1636 = {{2'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3633 = _T_3632 + _GEN_1636; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1637 = {{3'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3634 = _T_3633 + _GEN_1637; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1638 = {{4'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3635 = _T_3634 + _GEN_1638; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1639 = {{5'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3636 = _T_3635 + _GEN_1639; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1640 = {{6'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3637 = _T_3636 + _GEN_1640; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3638 = 8'h2 == _T_3637; // @[Conditional.scala 37:30]
  wire  _T_3640 = 8'h3 == _T_3637; // @[Conditional.scala 37:30]
  wire  _GEN_375 = _T_3638 ? regs[187] : _T_3640; // @[Conditional.scala 40:58]
  wire [1:0] _T_3649 = regs[171] + regs[172]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1641 = {{1'd0}, regs[173]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3650 = _T_3649 + _GEN_1641; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1642 = {{2'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3651 = _T_3650 + _GEN_1642; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1643 = {{3'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3652 = _T_3651 + _GEN_1643; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1644 = {{4'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3653 = _T_3652 + _GEN_1644; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1645 = {{5'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3654 = _T_3653 + _GEN_1645; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1646 = {{6'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3655 = _T_3654 + _GEN_1646; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3656 = 8'h2 == _T_3655; // @[Conditional.scala 37:30]
  wire  _T_3658 = 8'h3 == _T_3655; // @[Conditional.scala 37:30]
  wire  _GEN_377 = _T_3656 ? regs[188] : _T_3658; // @[Conditional.scala 40:58]
  wire [1:0] _T_3667 = regs[172] + regs[173]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1647 = {{1'd0}, regs[174]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3668 = _T_3667 + _GEN_1647; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1648 = {{2'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3669 = _T_3668 + _GEN_1648; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1649 = {{3'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3670 = _T_3669 + _GEN_1649; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1650 = {{4'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3671 = _T_3670 + _GEN_1650; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1651 = {{5'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3672 = _T_3671 + _GEN_1651; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1652 = {{6'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3673 = _T_3672 + _GEN_1652; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3674 = 8'h2 == _T_3673; // @[Conditional.scala 37:30]
  wire  _T_3676 = 8'h3 == _T_3673; // @[Conditional.scala 37:30]
  wire  _GEN_379 = _T_3674 ? regs[189] : _T_3676; // @[Conditional.scala 40:58]
  wire [1:0] _T_3685 = regs[173] + regs[174]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1653 = {{1'd0}, regs[175]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3686 = _T_3685 + _GEN_1653; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1654 = {{2'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3687 = _T_3686 + _GEN_1654; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1655 = {{3'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3688 = _T_3687 + _GEN_1655; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1656 = {{4'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3689 = _T_3688 + _GEN_1656; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1657 = {{5'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3690 = _T_3689 + _GEN_1657; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1658 = {{6'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3691 = _T_3690 + _GEN_1658; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3692 = 8'h2 == _T_3691; // @[Conditional.scala 37:30]
  wire  _T_3694 = 8'h3 == _T_3691; // @[Conditional.scala 37:30]
  wire  _GEN_381 = _T_3692 ? regs[190] : _T_3694; // @[Conditional.scala 40:58]
  wire [1:0] _T_3703 = regs[174] + regs[175]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1659 = {{1'd0}, regs[160]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3704 = _T_3703 + _GEN_1659; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1660 = {{2'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3705 = _T_3704 + _GEN_1660; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1661 = {{3'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3706 = _T_3705 + _GEN_1661; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1662 = {{4'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3707 = _T_3706 + _GEN_1662; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1663 = {{5'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3708 = _T_3707 + _GEN_1663; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1664 = {{6'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3709 = _T_3708 + _GEN_1664; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3710 = 8'h2 == _T_3709; // @[Conditional.scala 37:30]
  wire  _T_3712 = 8'h3 == _T_3709; // @[Conditional.scala 37:30]
  wire  _GEN_383 = _T_3710 ? regs[191] : _T_3712; // @[Conditional.scala 40:58]
  wire [1:0] _T_3721 = regs[191] + regs[176]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1665 = {{1'd0}, regs[177]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3722 = _T_3721 + _GEN_1665; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1666 = {{2'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3723 = _T_3722 + _GEN_1666; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1667 = {{3'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3724 = _T_3723 + _GEN_1667; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1668 = {{4'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3725 = _T_3724 + _GEN_1668; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1669 = {{5'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3726 = _T_3725 + _GEN_1669; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1670 = {{6'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3727 = _T_3726 + _GEN_1670; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3728 = 8'h2 == _T_3727; // @[Conditional.scala 37:30]
  wire  _T_3730 = 8'h3 == _T_3727; // @[Conditional.scala 37:30]
  wire  _GEN_385 = _T_3728 ? regs[192] : _T_3730; // @[Conditional.scala 40:58]
  wire [1:0] _T_3739 = regs[176] + regs[177]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1671 = {{1'd0}, regs[178]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3740 = _T_3739 + _GEN_1671; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1672 = {{2'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3741 = _T_3740 + _GEN_1672; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1673 = {{3'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3742 = _T_3741 + _GEN_1673; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1674 = {{4'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3743 = _T_3742 + _GEN_1674; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1675 = {{5'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3744 = _T_3743 + _GEN_1675; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1676 = {{6'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3745 = _T_3744 + _GEN_1676; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3746 = 8'h2 == _T_3745; // @[Conditional.scala 37:30]
  wire  _T_3748 = 8'h3 == _T_3745; // @[Conditional.scala 37:30]
  wire  _GEN_387 = _T_3746 ? regs[193] : _T_3748; // @[Conditional.scala 40:58]
  wire [1:0] _T_3757 = regs[177] + regs[178]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1677 = {{1'd0}, regs[179]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3758 = _T_3757 + _GEN_1677; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1678 = {{2'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3759 = _T_3758 + _GEN_1678; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1679 = {{3'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3760 = _T_3759 + _GEN_1679; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1680 = {{4'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3761 = _T_3760 + _GEN_1680; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1681 = {{5'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3762 = _T_3761 + _GEN_1681; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1682 = {{6'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3763 = _T_3762 + _GEN_1682; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3764 = 8'h2 == _T_3763; // @[Conditional.scala 37:30]
  wire  _T_3766 = 8'h3 == _T_3763; // @[Conditional.scala 37:30]
  wire  _GEN_389 = _T_3764 ? regs[194] : _T_3766; // @[Conditional.scala 40:58]
  wire [1:0] _T_3775 = regs[178] + regs[179]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1683 = {{1'd0}, regs[180]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3776 = _T_3775 + _GEN_1683; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1684 = {{2'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3777 = _T_3776 + _GEN_1684; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1685 = {{3'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3778 = _T_3777 + _GEN_1685; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1686 = {{4'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3779 = _T_3778 + _GEN_1686; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1687 = {{5'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3780 = _T_3779 + _GEN_1687; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1688 = {{6'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3781 = _T_3780 + _GEN_1688; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3782 = 8'h2 == _T_3781; // @[Conditional.scala 37:30]
  wire  _T_3784 = 8'h3 == _T_3781; // @[Conditional.scala 37:30]
  wire  _GEN_391 = _T_3782 ? regs[195] : _T_3784; // @[Conditional.scala 40:58]
  wire [1:0] _T_3793 = regs[179] + regs[180]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1689 = {{1'd0}, regs[181]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3794 = _T_3793 + _GEN_1689; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1690 = {{2'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3795 = _T_3794 + _GEN_1690; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1691 = {{3'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3796 = _T_3795 + _GEN_1691; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1692 = {{4'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3797 = _T_3796 + _GEN_1692; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1693 = {{5'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3798 = _T_3797 + _GEN_1693; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1694 = {{6'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3799 = _T_3798 + _GEN_1694; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3800 = 8'h2 == _T_3799; // @[Conditional.scala 37:30]
  wire  _T_3802 = 8'h3 == _T_3799; // @[Conditional.scala 37:30]
  wire  _GEN_393 = _T_3800 ? regs[196] : _T_3802; // @[Conditional.scala 40:58]
  wire [1:0] _T_3811 = regs[180] + regs[181]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1695 = {{1'd0}, regs[182]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3812 = _T_3811 + _GEN_1695; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1696 = {{2'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3813 = _T_3812 + _GEN_1696; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1697 = {{3'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3814 = _T_3813 + _GEN_1697; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1698 = {{4'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3815 = _T_3814 + _GEN_1698; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1699 = {{5'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3816 = _T_3815 + _GEN_1699; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1700 = {{6'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3817 = _T_3816 + _GEN_1700; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3818 = 8'h2 == _T_3817; // @[Conditional.scala 37:30]
  wire  _T_3820 = 8'h3 == _T_3817; // @[Conditional.scala 37:30]
  wire  _GEN_395 = _T_3818 ? regs[197] : _T_3820; // @[Conditional.scala 40:58]
  wire [1:0] _T_3829 = regs[181] + regs[182]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1701 = {{1'd0}, regs[183]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3830 = _T_3829 + _GEN_1701; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1702 = {{2'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3831 = _T_3830 + _GEN_1702; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1703 = {{3'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3832 = _T_3831 + _GEN_1703; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1704 = {{4'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3833 = _T_3832 + _GEN_1704; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1705 = {{5'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3834 = _T_3833 + _GEN_1705; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1706 = {{6'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3835 = _T_3834 + _GEN_1706; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3836 = 8'h2 == _T_3835; // @[Conditional.scala 37:30]
  wire  _T_3838 = 8'h3 == _T_3835; // @[Conditional.scala 37:30]
  wire  _GEN_397 = _T_3836 ? regs[198] : _T_3838; // @[Conditional.scala 40:58]
  wire [1:0] _T_3847 = regs[182] + regs[183]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1707 = {{1'd0}, regs[184]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3848 = _T_3847 + _GEN_1707; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1708 = {{2'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3849 = _T_3848 + _GEN_1708; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1709 = {{3'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3850 = _T_3849 + _GEN_1709; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1710 = {{4'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3851 = _T_3850 + _GEN_1710; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1711 = {{5'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3852 = _T_3851 + _GEN_1711; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1712 = {{6'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3853 = _T_3852 + _GEN_1712; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3854 = 8'h2 == _T_3853; // @[Conditional.scala 37:30]
  wire  _T_3856 = 8'h3 == _T_3853; // @[Conditional.scala 37:30]
  wire  _GEN_399 = _T_3854 ? regs[199] : _T_3856; // @[Conditional.scala 40:58]
  wire [1:0] _T_3865 = regs[183] + regs[184]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1713 = {{1'd0}, regs[185]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3866 = _T_3865 + _GEN_1713; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1714 = {{2'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3867 = _T_3866 + _GEN_1714; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1715 = {{3'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3868 = _T_3867 + _GEN_1715; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1716 = {{4'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3869 = _T_3868 + _GEN_1716; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1717 = {{5'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3870 = _T_3869 + _GEN_1717; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1718 = {{6'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3871 = _T_3870 + _GEN_1718; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3872 = 8'h2 == _T_3871; // @[Conditional.scala 37:30]
  wire  _T_3874 = 8'h3 == _T_3871; // @[Conditional.scala 37:30]
  wire  _GEN_401 = _T_3872 ? regs[200] : _T_3874; // @[Conditional.scala 40:58]
  wire [1:0] _T_3883 = regs[184] + regs[185]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1719 = {{1'd0}, regs[186]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3884 = _T_3883 + _GEN_1719; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1720 = {{2'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3885 = _T_3884 + _GEN_1720; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1721 = {{3'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3886 = _T_3885 + _GEN_1721; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1722 = {{4'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3887 = _T_3886 + _GEN_1722; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1723 = {{5'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3888 = _T_3887 + _GEN_1723; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1724 = {{6'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3889 = _T_3888 + _GEN_1724; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3890 = 8'h2 == _T_3889; // @[Conditional.scala 37:30]
  wire  _T_3892 = 8'h3 == _T_3889; // @[Conditional.scala 37:30]
  wire  _GEN_403 = _T_3890 ? regs[201] : _T_3892; // @[Conditional.scala 40:58]
  wire [1:0] _T_3901 = regs[185] + regs[186]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1725 = {{1'd0}, regs[187]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3902 = _T_3901 + _GEN_1725; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1726 = {{2'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3903 = _T_3902 + _GEN_1726; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1727 = {{3'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3904 = _T_3903 + _GEN_1727; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1728 = {{4'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3905 = _T_3904 + _GEN_1728; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1729 = {{5'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3906 = _T_3905 + _GEN_1729; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1730 = {{6'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3907 = _T_3906 + _GEN_1730; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3908 = 8'h2 == _T_3907; // @[Conditional.scala 37:30]
  wire  _T_3910 = 8'h3 == _T_3907; // @[Conditional.scala 37:30]
  wire  _GEN_405 = _T_3908 ? regs[202] : _T_3910; // @[Conditional.scala 40:58]
  wire [1:0] _T_3919 = regs[186] + regs[187]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1731 = {{1'd0}, regs[188]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3920 = _T_3919 + _GEN_1731; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1732 = {{2'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3921 = _T_3920 + _GEN_1732; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1733 = {{3'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3922 = _T_3921 + _GEN_1733; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1734 = {{4'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3923 = _T_3922 + _GEN_1734; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1735 = {{5'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3924 = _T_3923 + _GEN_1735; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1736 = {{6'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3925 = _T_3924 + _GEN_1736; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3926 = 8'h2 == _T_3925; // @[Conditional.scala 37:30]
  wire  _T_3928 = 8'h3 == _T_3925; // @[Conditional.scala 37:30]
  wire  _GEN_407 = _T_3926 ? regs[203] : _T_3928; // @[Conditional.scala 40:58]
  wire [1:0] _T_3937 = regs[187] + regs[188]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1737 = {{1'd0}, regs[189]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3938 = _T_3937 + _GEN_1737; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1738 = {{2'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3939 = _T_3938 + _GEN_1738; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1739 = {{3'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3940 = _T_3939 + _GEN_1739; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1740 = {{4'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3941 = _T_3940 + _GEN_1740; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1741 = {{5'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3942 = _T_3941 + _GEN_1741; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1742 = {{6'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3943 = _T_3942 + _GEN_1742; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3944 = 8'h2 == _T_3943; // @[Conditional.scala 37:30]
  wire  _T_3946 = 8'h3 == _T_3943; // @[Conditional.scala 37:30]
  wire  _GEN_409 = _T_3944 ? regs[204] : _T_3946; // @[Conditional.scala 40:58]
  wire [1:0] _T_3955 = regs[188] + regs[189]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1743 = {{1'd0}, regs[190]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3956 = _T_3955 + _GEN_1743; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1744 = {{2'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3957 = _T_3956 + _GEN_1744; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1745 = {{3'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3958 = _T_3957 + _GEN_1745; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1746 = {{4'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3959 = _T_3958 + _GEN_1746; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1747 = {{5'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3960 = _T_3959 + _GEN_1747; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1748 = {{6'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3961 = _T_3960 + _GEN_1748; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3962 = 8'h2 == _T_3961; // @[Conditional.scala 37:30]
  wire  _T_3964 = 8'h3 == _T_3961; // @[Conditional.scala 37:30]
  wire  _GEN_411 = _T_3962 ? regs[205] : _T_3964; // @[Conditional.scala 40:58]
  wire [1:0] _T_3973 = regs[189] + regs[190]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1749 = {{1'd0}, regs[191]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3974 = _T_3973 + _GEN_1749; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1750 = {{2'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3975 = _T_3974 + _GEN_1750; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1751 = {{3'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3976 = _T_3975 + _GEN_1751; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1752 = {{4'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3977 = _T_3976 + _GEN_1752; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1753 = {{5'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3978 = _T_3977 + _GEN_1753; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1754 = {{6'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3979 = _T_3978 + _GEN_1754; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3980 = 8'h2 == _T_3979; // @[Conditional.scala 37:30]
  wire  _T_3982 = 8'h3 == _T_3979; // @[Conditional.scala 37:30]
  wire  _GEN_413 = _T_3980 ? regs[206] : _T_3982; // @[Conditional.scala 40:58]
  wire [1:0] _T_3991 = regs[190] + regs[191]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1755 = {{1'd0}, regs[176]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_3992 = _T_3991 + _GEN_1755; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1756 = {{2'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_3993 = _T_3992 + _GEN_1756; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1757 = {{3'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_3994 = _T_3993 + _GEN_1757; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1758 = {{4'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_3995 = _T_3994 + _GEN_1758; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1759 = {{5'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_3996 = _T_3995 + _GEN_1759; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1760 = {{6'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_3997 = _T_3996 + _GEN_1760; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_3998 = 8'h2 == _T_3997; // @[Conditional.scala 37:30]
  wire  _T_4000 = 8'h3 == _T_3997; // @[Conditional.scala 37:30]
  wire  _GEN_415 = _T_3998 ? regs[207] : _T_4000; // @[Conditional.scala 40:58]
  wire [1:0] _T_4009 = regs[207] + regs[192]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1761 = {{1'd0}, regs[193]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4010 = _T_4009 + _GEN_1761; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1762 = {{2'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4011 = _T_4010 + _GEN_1762; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1763 = {{3'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4012 = _T_4011 + _GEN_1763; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1764 = {{4'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4013 = _T_4012 + _GEN_1764; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1765 = {{5'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4014 = _T_4013 + _GEN_1765; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1766 = {{6'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4015 = _T_4014 + _GEN_1766; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4016 = 8'h2 == _T_4015; // @[Conditional.scala 37:30]
  wire  _T_4018 = 8'h3 == _T_4015; // @[Conditional.scala 37:30]
  wire  _GEN_417 = _T_4016 ? regs[208] : _T_4018; // @[Conditional.scala 40:58]
  wire [1:0] _T_4027 = regs[192] + regs[193]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1767 = {{1'd0}, regs[194]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4028 = _T_4027 + _GEN_1767; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1768 = {{2'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4029 = _T_4028 + _GEN_1768; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1769 = {{3'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4030 = _T_4029 + _GEN_1769; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1770 = {{4'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4031 = _T_4030 + _GEN_1770; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1771 = {{5'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4032 = _T_4031 + _GEN_1771; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1772 = {{6'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4033 = _T_4032 + _GEN_1772; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4034 = 8'h2 == _T_4033; // @[Conditional.scala 37:30]
  wire  _T_4036 = 8'h3 == _T_4033; // @[Conditional.scala 37:30]
  wire  _GEN_419 = _T_4034 ? regs[209] : _T_4036; // @[Conditional.scala 40:58]
  wire [1:0] _T_4045 = regs[193] + regs[194]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1773 = {{1'd0}, regs[195]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4046 = _T_4045 + _GEN_1773; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1774 = {{2'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4047 = _T_4046 + _GEN_1774; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1775 = {{3'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4048 = _T_4047 + _GEN_1775; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1776 = {{4'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4049 = _T_4048 + _GEN_1776; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1777 = {{5'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4050 = _T_4049 + _GEN_1777; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1778 = {{6'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4051 = _T_4050 + _GEN_1778; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4052 = 8'h2 == _T_4051; // @[Conditional.scala 37:30]
  wire  _T_4054 = 8'h3 == _T_4051; // @[Conditional.scala 37:30]
  wire  _GEN_421 = _T_4052 ? regs[210] : _T_4054; // @[Conditional.scala 40:58]
  wire [1:0] _T_4063 = regs[194] + regs[195]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1779 = {{1'd0}, regs[196]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4064 = _T_4063 + _GEN_1779; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1780 = {{2'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4065 = _T_4064 + _GEN_1780; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1781 = {{3'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4066 = _T_4065 + _GEN_1781; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1782 = {{4'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4067 = _T_4066 + _GEN_1782; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1783 = {{5'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4068 = _T_4067 + _GEN_1783; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1784 = {{6'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4069 = _T_4068 + _GEN_1784; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4070 = 8'h2 == _T_4069; // @[Conditional.scala 37:30]
  wire  _T_4072 = 8'h3 == _T_4069; // @[Conditional.scala 37:30]
  wire  _GEN_423 = _T_4070 ? regs[211] : _T_4072; // @[Conditional.scala 40:58]
  wire [1:0] _T_4081 = regs[195] + regs[196]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1785 = {{1'd0}, regs[197]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4082 = _T_4081 + _GEN_1785; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1786 = {{2'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4083 = _T_4082 + _GEN_1786; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1787 = {{3'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4084 = _T_4083 + _GEN_1787; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1788 = {{4'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4085 = _T_4084 + _GEN_1788; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1789 = {{5'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4086 = _T_4085 + _GEN_1789; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1790 = {{6'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4087 = _T_4086 + _GEN_1790; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4088 = 8'h2 == _T_4087; // @[Conditional.scala 37:30]
  wire  _T_4090 = 8'h3 == _T_4087; // @[Conditional.scala 37:30]
  wire  _GEN_425 = _T_4088 ? regs[212] : _T_4090; // @[Conditional.scala 40:58]
  wire [1:0] _T_4099 = regs[196] + regs[197]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1791 = {{1'd0}, regs[198]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4100 = _T_4099 + _GEN_1791; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1792 = {{2'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4101 = _T_4100 + _GEN_1792; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1793 = {{3'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4102 = _T_4101 + _GEN_1793; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1794 = {{4'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4103 = _T_4102 + _GEN_1794; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1795 = {{5'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4104 = _T_4103 + _GEN_1795; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1796 = {{6'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4105 = _T_4104 + _GEN_1796; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4106 = 8'h2 == _T_4105; // @[Conditional.scala 37:30]
  wire  _T_4108 = 8'h3 == _T_4105; // @[Conditional.scala 37:30]
  wire  _GEN_427 = _T_4106 ? regs[213] : _T_4108; // @[Conditional.scala 40:58]
  wire [1:0] _T_4117 = regs[197] + regs[198]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1797 = {{1'd0}, regs[199]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4118 = _T_4117 + _GEN_1797; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1798 = {{2'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4119 = _T_4118 + _GEN_1798; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1799 = {{3'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4120 = _T_4119 + _GEN_1799; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1800 = {{4'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4121 = _T_4120 + _GEN_1800; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1801 = {{5'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4122 = _T_4121 + _GEN_1801; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1802 = {{6'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4123 = _T_4122 + _GEN_1802; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4124 = 8'h2 == _T_4123; // @[Conditional.scala 37:30]
  wire  _T_4126 = 8'h3 == _T_4123; // @[Conditional.scala 37:30]
  wire  _GEN_429 = _T_4124 ? regs[214] : _T_4126; // @[Conditional.scala 40:58]
  wire [1:0] _T_4135 = regs[198] + regs[199]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1803 = {{1'd0}, regs[200]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4136 = _T_4135 + _GEN_1803; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1804 = {{2'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4137 = _T_4136 + _GEN_1804; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1805 = {{3'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4138 = _T_4137 + _GEN_1805; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1806 = {{4'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4139 = _T_4138 + _GEN_1806; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1807 = {{5'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4140 = _T_4139 + _GEN_1807; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1808 = {{6'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4141 = _T_4140 + _GEN_1808; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4142 = 8'h2 == _T_4141; // @[Conditional.scala 37:30]
  wire  _T_4144 = 8'h3 == _T_4141; // @[Conditional.scala 37:30]
  wire  _GEN_431 = _T_4142 ? regs[215] : _T_4144; // @[Conditional.scala 40:58]
  wire [1:0] _T_4153 = regs[199] + regs[200]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1809 = {{1'd0}, regs[201]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4154 = _T_4153 + _GEN_1809; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1810 = {{2'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4155 = _T_4154 + _GEN_1810; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1811 = {{3'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4156 = _T_4155 + _GEN_1811; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1812 = {{4'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4157 = _T_4156 + _GEN_1812; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1813 = {{5'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4158 = _T_4157 + _GEN_1813; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1814 = {{6'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4159 = _T_4158 + _GEN_1814; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4160 = 8'h2 == _T_4159; // @[Conditional.scala 37:30]
  wire  _T_4162 = 8'h3 == _T_4159; // @[Conditional.scala 37:30]
  wire  _GEN_433 = _T_4160 ? regs[216] : _T_4162; // @[Conditional.scala 40:58]
  wire [1:0] _T_4171 = regs[200] + regs[201]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1815 = {{1'd0}, regs[202]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4172 = _T_4171 + _GEN_1815; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1816 = {{2'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4173 = _T_4172 + _GEN_1816; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1817 = {{3'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4174 = _T_4173 + _GEN_1817; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1818 = {{4'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4175 = _T_4174 + _GEN_1818; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1819 = {{5'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4176 = _T_4175 + _GEN_1819; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1820 = {{6'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4177 = _T_4176 + _GEN_1820; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4178 = 8'h2 == _T_4177; // @[Conditional.scala 37:30]
  wire  _T_4180 = 8'h3 == _T_4177; // @[Conditional.scala 37:30]
  wire  _GEN_435 = _T_4178 ? regs[217] : _T_4180; // @[Conditional.scala 40:58]
  wire [1:0] _T_4189 = regs[201] + regs[202]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1821 = {{1'd0}, regs[203]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4190 = _T_4189 + _GEN_1821; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1822 = {{2'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4191 = _T_4190 + _GEN_1822; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1823 = {{3'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4192 = _T_4191 + _GEN_1823; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1824 = {{4'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4193 = _T_4192 + _GEN_1824; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1825 = {{5'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4194 = _T_4193 + _GEN_1825; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1826 = {{6'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4195 = _T_4194 + _GEN_1826; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4196 = 8'h2 == _T_4195; // @[Conditional.scala 37:30]
  wire  _T_4198 = 8'h3 == _T_4195; // @[Conditional.scala 37:30]
  wire  _GEN_437 = _T_4196 ? regs[218] : _T_4198; // @[Conditional.scala 40:58]
  wire [1:0] _T_4207 = regs[202] + regs[203]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1827 = {{1'd0}, regs[204]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4208 = _T_4207 + _GEN_1827; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1828 = {{2'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4209 = _T_4208 + _GEN_1828; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1829 = {{3'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4210 = _T_4209 + _GEN_1829; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1830 = {{4'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4211 = _T_4210 + _GEN_1830; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1831 = {{5'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4212 = _T_4211 + _GEN_1831; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1832 = {{6'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4213 = _T_4212 + _GEN_1832; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4214 = 8'h2 == _T_4213; // @[Conditional.scala 37:30]
  wire  _T_4216 = 8'h3 == _T_4213; // @[Conditional.scala 37:30]
  wire  _GEN_439 = _T_4214 ? regs[219] : _T_4216; // @[Conditional.scala 40:58]
  wire [1:0] _T_4225 = regs[203] + regs[204]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1833 = {{1'd0}, regs[205]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4226 = _T_4225 + _GEN_1833; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1834 = {{2'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4227 = _T_4226 + _GEN_1834; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1835 = {{3'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4228 = _T_4227 + _GEN_1835; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1836 = {{4'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4229 = _T_4228 + _GEN_1836; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1837 = {{5'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4230 = _T_4229 + _GEN_1837; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1838 = {{6'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4231 = _T_4230 + _GEN_1838; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4232 = 8'h2 == _T_4231; // @[Conditional.scala 37:30]
  wire  _T_4234 = 8'h3 == _T_4231; // @[Conditional.scala 37:30]
  wire  _GEN_441 = _T_4232 ? regs[220] : _T_4234; // @[Conditional.scala 40:58]
  wire [1:0] _T_4243 = regs[204] + regs[205]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1839 = {{1'd0}, regs[206]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4244 = _T_4243 + _GEN_1839; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1840 = {{2'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4245 = _T_4244 + _GEN_1840; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1841 = {{3'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4246 = _T_4245 + _GEN_1841; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1842 = {{4'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4247 = _T_4246 + _GEN_1842; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1843 = {{5'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4248 = _T_4247 + _GEN_1843; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1844 = {{6'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4249 = _T_4248 + _GEN_1844; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4250 = 8'h2 == _T_4249; // @[Conditional.scala 37:30]
  wire  _T_4252 = 8'h3 == _T_4249; // @[Conditional.scala 37:30]
  wire  _GEN_443 = _T_4250 ? regs[221] : _T_4252; // @[Conditional.scala 40:58]
  wire [1:0] _T_4261 = regs[205] + regs[206]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1845 = {{1'd0}, regs[207]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4262 = _T_4261 + _GEN_1845; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1846 = {{2'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4263 = _T_4262 + _GEN_1846; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1847 = {{3'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4264 = _T_4263 + _GEN_1847; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1848 = {{4'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4265 = _T_4264 + _GEN_1848; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1849 = {{5'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4266 = _T_4265 + _GEN_1849; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1850 = {{6'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4267 = _T_4266 + _GEN_1850; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4268 = 8'h2 == _T_4267; // @[Conditional.scala 37:30]
  wire  _T_4270 = 8'h3 == _T_4267; // @[Conditional.scala 37:30]
  wire  _GEN_445 = _T_4268 ? regs[222] : _T_4270; // @[Conditional.scala 40:58]
  wire [1:0] _T_4279 = regs[206] + regs[207]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1851 = {{1'd0}, regs[192]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4280 = _T_4279 + _GEN_1851; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1852 = {{2'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4281 = _T_4280 + _GEN_1852; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1853 = {{3'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4282 = _T_4281 + _GEN_1853; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1854 = {{4'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4283 = _T_4282 + _GEN_1854; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1855 = {{5'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4284 = _T_4283 + _GEN_1855; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1856 = {{6'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4285 = _T_4284 + _GEN_1856; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4286 = 8'h2 == _T_4285; // @[Conditional.scala 37:30]
  wire  _T_4288 = 8'h3 == _T_4285; // @[Conditional.scala 37:30]
  wire  _GEN_447 = _T_4286 ? regs[223] : _T_4288; // @[Conditional.scala 40:58]
  wire [1:0] _T_4297 = regs[223] + regs[208]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1857 = {{1'd0}, regs[209]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4298 = _T_4297 + _GEN_1857; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1858 = {{2'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4299 = _T_4298 + _GEN_1858; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1859 = {{3'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4300 = _T_4299 + _GEN_1859; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1860 = {{4'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4301 = _T_4300 + _GEN_1860; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1861 = {{5'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4302 = _T_4301 + _GEN_1861; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1862 = {{6'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4303 = _T_4302 + _GEN_1862; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4304 = 8'h2 == _T_4303; // @[Conditional.scala 37:30]
  wire  _T_4306 = 8'h3 == _T_4303; // @[Conditional.scala 37:30]
  wire  _GEN_449 = _T_4304 ? regs[224] : _T_4306; // @[Conditional.scala 40:58]
  wire [1:0] _T_4315 = regs[208] + regs[209]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1863 = {{1'd0}, regs[210]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4316 = _T_4315 + _GEN_1863; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1864 = {{2'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4317 = _T_4316 + _GEN_1864; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1865 = {{3'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4318 = _T_4317 + _GEN_1865; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1866 = {{4'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4319 = _T_4318 + _GEN_1866; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1867 = {{5'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4320 = _T_4319 + _GEN_1867; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1868 = {{6'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4321 = _T_4320 + _GEN_1868; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4322 = 8'h2 == _T_4321; // @[Conditional.scala 37:30]
  wire  _T_4324 = 8'h3 == _T_4321; // @[Conditional.scala 37:30]
  wire  _GEN_451 = _T_4322 ? regs[225] : _T_4324; // @[Conditional.scala 40:58]
  wire [1:0] _T_4333 = regs[209] + regs[210]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1869 = {{1'd0}, regs[211]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4334 = _T_4333 + _GEN_1869; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1870 = {{2'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4335 = _T_4334 + _GEN_1870; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1871 = {{3'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4336 = _T_4335 + _GEN_1871; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1872 = {{4'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4337 = _T_4336 + _GEN_1872; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1873 = {{5'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4338 = _T_4337 + _GEN_1873; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1874 = {{6'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4339 = _T_4338 + _GEN_1874; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4340 = 8'h2 == _T_4339; // @[Conditional.scala 37:30]
  wire  _T_4342 = 8'h3 == _T_4339; // @[Conditional.scala 37:30]
  wire  _GEN_453 = _T_4340 ? regs[226] : _T_4342; // @[Conditional.scala 40:58]
  wire [1:0] _T_4351 = regs[210] + regs[211]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1875 = {{1'd0}, regs[212]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4352 = _T_4351 + _GEN_1875; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1876 = {{2'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4353 = _T_4352 + _GEN_1876; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1877 = {{3'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4354 = _T_4353 + _GEN_1877; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1878 = {{4'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4355 = _T_4354 + _GEN_1878; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1879 = {{5'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4356 = _T_4355 + _GEN_1879; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1880 = {{6'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4357 = _T_4356 + _GEN_1880; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4358 = 8'h2 == _T_4357; // @[Conditional.scala 37:30]
  wire  _T_4360 = 8'h3 == _T_4357; // @[Conditional.scala 37:30]
  wire  _GEN_455 = _T_4358 ? regs[227] : _T_4360; // @[Conditional.scala 40:58]
  wire [1:0] _T_4369 = regs[211] + regs[212]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1881 = {{1'd0}, regs[213]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4370 = _T_4369 + _GEN_1881; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1882 = {{2'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4371 = _T_4370 + _GEN_1882; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1883 = {{3'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4372 = _T_4371 + _GEN_1883; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1884 = {{4'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4373 = _T_4372 + _GEN_1884; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1885 = {{5'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4374 = _T_4373 + _GEN_1885; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1886 = {{6'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4375 = _T_4374 + _GEN_1886; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4376 = 8'h2 == _T_4375; // @[Conditional.scala 37:30]
  wire  _T_4378 = 8'h3 == _T_4375; // @[Conditional.scala 37:30]
  wire  _GEN_457 = _T_4376 ? regs[228] : _T_4378; // @[Conditional.scala 40:58]
  wire [1:0] _T_4387 = regs[212] + regs[213]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1887 = {{1'd0}, regs[214]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4388 = _T_4387 + _GEN_1887; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1888 = {{2'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4389 = _T_4388 + _GEN_1888; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1889 = {{3'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4390 = _T_4389 + _GEN_1889; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1890 = {{4'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4391 = _T_4390 + _GEN_1890; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1891 = {{5'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4392 = _T_4391 + _GEN_1891; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1892 = {{6'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4393 = _T_4392 + _GEN_1892; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4394 = 8'h2 == _T_4393; // @[Conditional.scala 37:30]
  wire  _T_4396 = 8'h3 == _T_4393; // @[Conditional.scala 37:30]
  wire  _GEN_459 = _T_4394 ? regs[229] : _T_4396; // @[Conditional.scala 40:58]
  wire [1:0] _T_4405 = regs[213] + regs[214]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1893 = {{1'd0}, regs[215]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4406 = _T_4405 + _GEN_1893; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1894 = {{2'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4407 = _T_4406 + _GEN_1894; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1895 = {{3'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4408 = _T_4407 + _GEN_1895; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1896 = {{4'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4409 = _T_4408 + _GEN_1896; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1897 = {{5'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4410 = _T_4409 + _GEN_1897; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1898 = {{6'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4411 = _T_4410 + _GEN_1898; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4412 = 8'h2 == _T_4411; // @[Conditional.scala 37:30]
  wire  _T_4414 = 8'h3 == _T_4411; // @[Conditional.scala 37:30]
  wire  _GEN_461 = _T_4412 ? regs[230] : _T_4414; // @[Conditional.scala 40:58]
  wire [1:0] _T_4423 = regs[214] + regs[215]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1899 = {{1'd0}, regs[216]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4424 = _T_4423 + _GEN_1899; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1900 = {{2'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4425 = _T_4424 + _GEN_1900; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1901 = {{3'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4426 = _T_4425 + _GEN_1901; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1902 = {{4'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4427 = _T_4426 + _GEN_1902; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1903 = {{5'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4428 = _T_4427 + _GEN_1903; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1904 = {{6'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4429 = _T_4428 + _GEN_1904; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4430 = 8'h2 == _T_4429; // @[Conditional.scala 37:30]
  wire  _T_4432 = 8'h3 == _T_4429; // @[Conditional.scala 37:30]
  wire  _GEN_463 = _T_4430 ? regs[231] : _T_4432; // @[Conditional.scala 40:58]
  wire [1:0] _T_4441 = regs[215] + regs[216]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1905 = {{1'd0}, regs[217]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4442 = _T_4441 + _GEN_1905; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1906 = {{2'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4443 = _T_4442 + _GEN_1906; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1907 = {{3'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4444 = _T_4443 + _GEN_1907; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1908 = {{4'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4445 = _T_4444 + _GEN_1908; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1909 = {{5'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4446 = _T_4445 + _GEN_1909; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1910 = {{6'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4447 = _T_4446 + _GEN_1910; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4448 = 8'h2 == _T_4447; // @[Conditional.scala 37:30]
  wire  _T_4450 = 8'h3 == _T_4447; // @[Conditional.scala 37:30]
  wire  _GEN_465 = _T_4448 ? regs[232] : _T_4450; // @[Conditional.scala 40:58]
  wire [1:0] _T_4459 = regs[216] + regs[217]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1911 = {{1'd0}, regs[218]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4460 = _T_4459 + _GEN_1911; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1912 = {{2'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4461 = _T_4460 + _GEN_1912; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1913 = {{3'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4462 = _T_4461 + _GEN_1913; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1914 = {{4'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4463 = _T_4462 + _GEN_1914; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1915 = {{5'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4464 = _T_4463 + _GEN_1915; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1916 = {{6'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4465 = _T_4464 + _GEN_1916; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4466 = 8'h2 == _T_4465; // @[Conditional.scala 37:30]
  wire  _T_4468 = 8'h3 == _T_4465; // @[Conditional.scala 37:30]
  wire  _GEN_467 = _T_4466 ? regs[233] : _T_4468; // @[Conditional.scala 40:58]
  wire [1:0] _T_4477 = regs[217] + regs[218]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1917 = {{1'd0}, regs[219]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4478 = _T_4477 + _GEN_1917; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1918 = {{2'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4479 = _T_4478 + _GEN_1918; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1919 = {{3'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4480 = _T_4479 + _GEN_1919; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1920 = {{4'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4481 = _T_4480 + _GEN_1920; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1921 = {{5'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4482 = _T_4481 + _GEN_1921; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1922 = {{6'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4483 = _T_4482 + _GEN_1922; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4484 = 8'h2 == _T_4483; // @[Conditional.scala 37:30]
  wire  _T_4486 = 8'h3 == _T_4483; // @[Conditional.scala 37:30]
  wire  _GEN_469 = _T_4484 ? regs[234] : _T_4486; // @[Conditional.scala 40:58]
  wire [1:0] _T_4495 = regs[218] + regs[219]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1923 = {{1'd0}, regs[220]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4496 = _T_4495 + _GEN_1923; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1924 = {{2'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4497 = _T_4496 + _GEN_1924; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1925 = {{3'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4498 = _T_4497 + _GEN_1925; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1926 = {{4'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4499 = _T_4498 + _GEN_1926; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1927 = {{5'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4500 = _T_4499 + _GEN_1927; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1928 = {{6'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4501 = _T_4500 + _GEN_1928; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4502 = 8'h2 == _T_4501; // @[Conditional.scala 37:30]
  wire  _T_4504 = 8'h3 == _T_4501; // @[Conditional.scala 37:30]
  wire  _GEN_471 = _T_4502 ? regs[235] : _T_4504; // @[Conditional.scala 40:58]
  wire [1:0] _T_4513 = regs[219] + regs[220]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1929 = {{1'd0}, regs[221]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4514 = _T_4513 + _GEN_1929; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1930 = {{2'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4515 = _T_4514 + _GEN_1930; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1931 = {{3'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4516 = _T_4515 + _GEN_1931; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1932 = {{4'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4517 = _T_4516 + _GEN_1932; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1933 = {{5'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4518 = _T_4517 + _GEN_1933; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1934 = {{6'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4519 = _T_4518 + _GEN_1934; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4520 = 8'h2 == _T_4519; // @[Conditional.scala 37:30]
  wire  _T_4522 = 8'h3 == _T_4519; // @[Conditional.scala 37:30]
  wire  _GEN_473 = _T_4520 ? regs[236] : _T_4522; // @[Conditional.scala 40:58]
  wire [1:0] _T_4531 = regs[220] + regs[221]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1935 = {{1'd0}, regs[222]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4532 = _T_4531 + _GEN_1935; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1936 = {{2'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4533 = _T_4532 + _GEN_1936; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1937 = {{3'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4534 = _T_4533 + _GEN_1937; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1938 = {{4'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4535 = _T_4534 + _GEN_1938; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1939 = {{5'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4536 = _T_4535 + _GEN_1939; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1940 = {{6'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4537 = _T_4536 + _GEN_1940; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4538 = 8'h2 == _T_4537; // @[Conditional.scala 37:30]
  wire  _T_4540 = 8'h3 == _T_4537; // @[Conditional.scala 37:30]
  wire  _GEN_475 = _T_4538 ? regs[237] : _T_4540; // @[Conditional.scala 40:58]
  wire [1:0] _T_4549 = regs[221] + regs[222]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1941 = {{1'd0}, regs[223]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4550 = _T_4549 + _GEN_1941; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1942 = {{2'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4551 = _T_4550 + _GEN_1942; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1943 = {{3'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4552 = _T_4551 + _GEN_1943; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1944 = {{4'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4553 = _T_4552 + _GEN_1944; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1945 = {{5'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4554 = _T_4553 + _GEN_1945; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1946 = {{6'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4555 = _T_4554 + _GEN_1946; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4556 = 8'h2 == _T_4555; // @[Conditional.scala 37:30]
  wire  _T_4558 = 8'h3 == _T_4555; // @[Conditional.scala 37:30]
  wire  _GEN_477 = _T_4556 ? regs[238] : _T_4558; // @[Conditional.scala 40:58]
  wire [1:0] _T_4567 = regs[222] + regs[223]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1947 = {{1'd0}, regs[208]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4568 = _T_4567 + _GEN_1947; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1948 = {{2'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4569 = _T_4568 + _GEN_1948; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1949 = {{3'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4570 = _T_4569 + _GEN_1949; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1950 = {{4'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4571 = _T_4570 + _GEN_1950; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1951 = {{5'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4572 = _T_4571 + _GEN_1951; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1952 = {{6'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4573 = _T_4572 + _GEN_1952; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4574 = 8'h2 == _T_4573; // @[Conditional.scala 37:30]
  wire  _T_4576 = 8'h3 == _T_4573; // @[Conditional.scala 37:30]
  wire  _GEN_479 = _T_4574 ? regs[239] : _T_4576; // @[Conditional.scala 40:58]
  wire [1:0] _T_4585 = regs[239] + regs[224]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1953 = {{1'd0}, regs[225]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4586 = _T_4585 + _GEN_1953; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1954 = {{2'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4587 = _T_4586 + _GEN_1954; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1955 = {{3'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4588 = _T_4587 + _GEN_1955; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1956 = {{4'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4589 = _T_4588 + _GEN_1956; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1957 = {{5'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4590 = _T_4589 + _GEN_1957; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1958 = {{6'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4591 = _T_4590 + _GEN_1958; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4592 = 8'h2 == _T_4591; // @[Conditional.scala 37:30]
  wire  _T_4594 = 8'h3 == _T_4591; // @[Conditional.scala 37:30]
  wire  _GEN_481 = _T_4592 ? regs[240] : _T_4594; // @[Conditional.scala 40:58]
  wire [1:0] _T_4603 = regs[224] + regs[225]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1959 = {{1'd0}, regs[226]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4604 = _T_4603 + _GEN_1959; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1960 = {{2'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4605 = _T_4604 + _GEN_1960; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1961 = {{3'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4606 = _T_4605 + _GEN_1961; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1962 = {{4'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4607 = _T_4606 + _GEN_1962; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1963 = {{5'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4608 = _T_4607 + _GEN_1963; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1964 = {{6'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4609 = _T_4608 + _GEN_1964; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4610 = 8'h2 == _T_4609; // @[Conditional.scala 37:30]
  wire  _T_4612 = 8'h3 == _T_4609; // @[Conditional.scala 37:30]
  wire  _GEN_483 = _T_4610 ? regs[241] : _T_4612; // @[Conditional.scala 40:58]
  wire [1:0] _T_4621 = regs[225] + regs[226]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1965 = {{1'd0}, regs[227]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4622 = _T_4621 + _GEN_1965; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1966 = {{2'd0}, regs[241]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4623 = _T_4622 + _GEN_1966; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1967 = {{3'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4624 = _T_4623 + _GEN_1967; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1968 = {{4'd0}, regs[1]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4625 = _T_4624 + _GEN_1968; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1969 = {{5'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4626 = _T_4625 + _GEN_1969; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1970 = {{6'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4627 = _T_4626 + _GEN_1970; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4628 = 8'h2 == _T_4627; // @[Conditional.scala 37:30]
  wire  _T_4630 = 8'h3 == _T_4627; // @[Conditional.scala 37:30]
  wire  _GEN_485 = _T_4628 ? regs[242] : _T_4630; // @[Conditional.scala 40:58]
  wire [1:0] _T_4639 = regs[226] + regs[227]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1971 = {{1'd0}, regs[228]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4640 = _T_4639 + _GEN_1971; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1972 = {{2'd0}, regs[242]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4641 = _T_4640 + _GEN_1972; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1973 = {{3'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4642 = _T_4641 + _GEN_1973; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1974 = {{4'd0}, regs[2]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4643 = _T_4642 + _GEN_1974; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1975 = {{5'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4644 = _T_4643 + _GEN_1975; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1976 = {{6'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4645 = _T_4644 + _GEN_1976; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4646 = 8'h2 == _T_4645; // @[Conditional.scala 37:30]
  wire  _T_4648 = 8'h3 == _T_4645; // @[Conditional.scala 37:30]
  wire  _GEN_487 = _T_4646 ? regs[243] : _T_4648; // @[Conditional.scala 40:58]
  wire [1:0] _T_4657 = regs[227] + regs[228]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1977 = {{1'd0}, regs[229]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4658 = _T_4657 + _GEN_1977; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1978 = {{2'd0}, regs[243]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4659 = _T_4658 + _GEN_1978; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1979 = {{3'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4660 = _T_4659 + _GEN_1979; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1980 = {{4'd0}, regs[3]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4661 = _T_4660 + _GEN_1980; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1981 = {{5'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4662 = _T_4661 + _GEN_1981; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1982 = {{6'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4663 = _T_4662 + _GEN_1982; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4664 = 8'h2 == _T_4663; // @[Conditional.scala 37:30]
  wire  _T_4666 = 8'h3 == _T_4663; // @[Conditional.scala 37:30]
  wire  _GEN_489 = _T_4664 ? regs[244] : _T_4666; // @[Conditional.scala 40:58]
  wire [1:0] _T_4675 = regs[228] + regs[229]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1983 = {{1'd0}, regs[230]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4676 = _T_4675 + _GEN_1983; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1984 = {{2'd0}, regs[244]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4677 = _T_4676 + _GEN_1984; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1985 = {{3'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4678 = _T_4677 + _GEN_1985; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1986 = {{4'd0}, regs[4]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4679 = _T_4678 + _GEN_1986; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1987 = {{5'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4680 = _T_4679 + _GEN_1987; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1988 = {{6'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4681 = _T_4680 + _GEN_1988; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4682 = 8'h2 == _T_4681; // @[Conditional.scala 37:30]
  wire  _T_4684 = 8'h3 == _T_4681; // @[Conditional.scala 37:30]
  wire  _GEN_491 = _T_4682 ? regs[245] : _T_4684; // @[Conditional.scala 40:58]
  wire [1:0] _T_4693 = regs[229] + regs[230]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1989 = {{1'd0}, regs[231]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4694 = _T_4693 + _GEN_1989; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1990 = {{2'd0}, regs[245]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4695 = _T_4694 + _GEN_1990; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1991 = {{3'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4696 = _T_4695 + _GEN_1991; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1992 = {{4'd0}, regs[5]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4697 = _T_4696 + _GEN_1992; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1993 = {{5'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4698 = _T_4697 + _GEN_1993; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_1994 = {{6'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4699 = _T_4698 + _GEN_1994; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4700 = 8'h2 == _T_4699; // @[Conditional.scala 37:30]
  wire  _T_4702 = 8'h3 == _T_4699; // @[Conditional.scala 37:30]
  wire  _GEN_493 = _T_4700 ? regs[246] : _T_4702; // @[Conditional.scala 40:58]
  wire [1:0] _T_4711 = regs[230] + regs[231]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_1995 = {{1'd0}, regs[232]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4712 = _T_4711 + _GEN_1995; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_1996 = {{2'd0}, regs[246]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4713 = _T_4712 + _GEN_1996; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_1997 = {{3'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4714 = _T_4713 + _GEN_1997; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_1998 = {{4'd0}, regs[6]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4715 = _T_4714 + _GEN_1998; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_1999 = {{5'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4716 = _T_4715 + _GEN_1999; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2000 = {{6'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4717 = _T_4716 + _GEN_2000; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4718 = 8'h2 == _T_4717; // @[Conditional.scala 37:30]
  wire  _T_4720 = 8'h3 == _T_4717; // @[Conditional.scala 37:30]
  wire  _GEN_495 = _T_4718 ? regs[247] : _T_4720; // @[Conditional.scala 40:58]
  wire [1:0] _T_4729 = regs[231] + regs[232]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2001 = {{1'd0}, regs[233]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4730 = _T_4729 + _GEN_2001; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2002 = {{2'd0}, regs[247]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4731 = _T_4730 + _GEN_2002; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2003 = {{3'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4732 = _T_4731 + _GEN_2003; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2004 = {{4'd0}, regs[7]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4733 = _T_4732 + _GEN_2004; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2005 = {{5'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4734 = _T_4733 + _GEN_2005; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2006 = {{6'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4735 = _T_4734 + _GEN_2006; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4736 = 8'h2 == _T_4735; // @[Conditional.scala 37:30]
  wire  _T_4738 = 8'h3 == _T_4735; // @[Conditional.scala 37:30]
  wire  _GEN_497 = _T_4736 ? regs[248] : _T_4738; // @[Conditional.scala 40:58]
  wire [1:0] _T_4747 = regs[232] + regs[233]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2007 = {{1'd0}, regs[234]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4748 = _T_4747 + _GEN_2007; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2008 = {{2'd0}, regs[248]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4749 = _T_4748 + _GEN_2008; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2009 = {{3'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4750 = _T_4749 + _GEN_2009; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2010 = {{4'd0}, regs[8]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4751 = _T_4750 + _GEN_2010; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2011 = {{5'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4752 = _T_4751 + _GEN_2011; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2012 = {{6'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4753 = _T_4752 + _GEN_2012; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4754 = 8'h2 == _T_4753; // @[Conditional.scala 37:30]
  wire  _T_4756 = 8'h3 == _T_4753; // @[Conditional.scala 37:30]
  wire  _GEN_499 = _T_4754 ? regs[249] : _T_4756; // @[Conditional.scala 40:58]
  wire [1:0] _T_4765 = regs[233] + regs[234]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2013 = {{1'd0}, regs[235]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4766 = _T_4765 + _GEN_2013; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2014 = {{2'd0}, regs[249]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4767 = _T_4766 + _GEN_2014; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2015 = {{3'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4768 = _T_4767 + _GEN_2015; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2016 = {{4'd0}, regs[9]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4769 = _T_4768 + _GEN_2016; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2017 = {{5'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4770 = _T_4769 + _GEN_2017; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2018 = {{6'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4771 = _T_4770 + _GEN_2018; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4772 = 8'h2 == _T_4771; // @[Conditional.scala 37:30]
  wire  _T_4774 = 8'h3 == _T_4771; // @[Conditional.scala 37:30]
  wire  _GEN_501 = _T_4772 ? regs[250] : _T_4774; // @[Conditional.scala 40:58]
  wire [1:0] _T_4783 = regs[234] + regs[235]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2019 = {{1'd0}, regs[236]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4784 = _T_4783 + _GEN_2019; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2020 = {{2'd0}, regs[250]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4785 = _T_4784 + _GEN_2020; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2021 = {{3'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4786 = _T_4785 + _GEN_2021; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2022 = {{4'd0}, regs[10]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4787 = _T_4786 + _GEN_2022; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2023 = {{5'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4788 = _T_4787 + _GEN_2023; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2024 = {{6'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4789 = _T_4788 + _GEN_2024; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4790 = 8'h2 == _T_4789; // @[Conditional.scala 37:30]
  wire  _T_4792 = 8'h3 == _T_4789; // @[Conditional.scala 37:30]
  wire  _GEN_503 = _T_4790 ? regs[251] : _T_4792; // @[Conditional.scala 40:58]
  wire [1:0] _T_4801 = regs[235] + regs[236]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2025 = {{1'd0}, regs[237]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4802 = _T_4801 + _GEN_2025; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2026 = {{2'd0}, regs[251]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4803 = _T_4802 + _GEN_2026; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2027 = {{3'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4804 = _T_4803 + _GEN_2027; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2028 = {{4'd0}, regs[11]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4805 = _T_4804 + _GEN_2028; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2029 = {{5'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4806 = _T_4805 + _GEN_2029; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2030 = {{6'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4807 = _T_4806 + _GEN_2030; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4808 = 8'h2 == _T_4807; // @[Conditional.scala 37:30]
  wire  _T_4810 = 8'h3 == _T_4807; // @[Conditional.scala 37:30]
  wire  _GEN_505 = _T_4808 ? regs[252] : _T_4810; // @[Conditional.scala 40:58]
  wire [1:0] _T_4819 = regs[236] + regs[237]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2031 = {{1'd0}, regs[238]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4820 = _T_4819 + _GEN_2031; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2032 = {{2'd0}, regs[252]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4821 = _T_4820 + _GEN_2032; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2033 = {{3'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4822 = _T_4821 + _GEN_2033; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2034 = {{4'd0}, regs[12]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4823 = _T_4822 + _GEN_2034; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2035 = {{5'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4824 = _T_4823 + _GEN_2035; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2036 = {{6'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4825 = _T_4824 + _GEN_2036; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4826 = 8'h2 == _T_4825; // @[Conditional.scala 37:30]
  wire  _T_4828 = 8'h3 == _T_4825; // @[Conditional.scala 37:30]
  wire  _GEN_507 = _T_4826 ? regs[253] : _T_4828; // @[Conditional.scala 40:58]
  wire [1:0] _T_4837 = regs[237] + regs[238]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2037 = {{1'd0}, regs[239]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4838 = _T_4837 + _GEN_2037; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2038 = {{2'd0}, regs[253]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4839 = _T_4838 + _GEN_2038; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2039 = {{3'd0}, regs[255]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4840 = _T_4839 + _GEN_2039; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2040 = {{4'd0}, regs[13]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4841 = _T_4840 + _GEN_2040; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2041 = {{5'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4842 = _T_4841 + _GEN_2041; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2042 = {{6'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4843 = _T_4842 + _GEN_2042; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4844 = 8'h2 == _T_4843; // @[Conditional.scala 37:30]
  wire  _T_4846 = 8'h3 == _T_4843; // @[Conditional.scala 37:30]
  wire  _GEN_509 = _T_4844 ? regs[254] : _T_4846; // @[Conditional.scala 40:58]
  wire [1:0] _T_4855 = regs[238] + regs[239]; // @[ConwaylifeBetter.scala 29:21]
  wire [1:0] _GEN_2043 = {{1'd0}, regs[224]}; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _T_4856 = _T_4855 + _GEN_2043; // @[ConwaylifeBetter.scala 29:21]
  wire [2:0] _GEN_2044 = {{2'd0}, regs[254]}; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _T_4857 = _T_4856 + _GEN_2044; // @[ConwaylifeBetter.scala 29:21]
  wire [3:0] _GEN_2045 = {{3'd0}, regs[240]}; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _T_4858 = _T_4857 + _GEN_2045; // @[ConwaylifeBetter.scala 29:21]
  wire [4:0] _GEN_2046 = {{4'd0}, regs[14]}; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _T_4859 = _T_4858 + _GEN_2046; // @[ConwaylifeBetter.scala 29:21]
  wire [5:0] _GEN_2047 = {{5'd0}, regs[15]}; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _T_4860 = _T_4859 + _GEN_2047; // @[ConwaylifeBetter.scala 29:21]
  wire [6:0] _GEN_2048 = {{6'd0}, regs[0]}; // @[ConwaylifeBetter.scala 29:21]
  wire [7:0] _T_4861 = _T_4860 + _GEN_2048; // @[ConwaylifeBetter.scala 29:21]
  wire  _T_4862 = 8'h2 == _T_4861; // @[Conditional.scala 37:30]
  wire  _T_4864 = 8'h3 == _T_4861; // @[Conditional.scala 37:30]
  wire  _GEN_511 = _T_4862 ? regs[255] : _T_4864; // @[Conditional.scala 40:58]
  wire [7:0] _T_4871 = {_GEN_15,_GEN_13,_GEN_11,_GEN_9,_GEN_7,_GEN_5,_GEN_3,_GEN_1}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_4879 = {_GEN_31,_GEN_29,_GEN_27,_GEN_25,_GEN_23,_GEN_21,_GEN_19,_GEN_17,_T_4871}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4886 = {_GEN_47,_GEN_45,_GEN_43,_GEN_41,_GEN_39,_GEN_37,_GEN_35,_GEN_33}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_4895 = {_GEN_63,_GEN_61,_GEN_59,_GEN_57,_GEN_55,_GEN_53,_GEN_51,_GEN_49,_T_4886,_T_4879}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4902 = {_GEN_79,_GEN_77,_GEN_75,_GEN_73,_GEN_71,_GEN_69,_GEN_67,_GEN_65}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_4910 = {_GEN_95,_GEN_93,_GEN_91,_GEN_89,_GEN_87,_GEN_85,_GEN_83,_GEN_81,_T_4902}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4917 = {_GEN_111,_GEN_109,_GEN_107,_GEN_105,_GEN_103,_GEN_101,_GEN_99,_GEN_97}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_4926 = {_GEN_127,_GEN_125,_GEN_123,_GEN_121,_GEN_119,_GEN_117,_GEN_115,_GEN_113,_T_4917,_T_4910}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4934 = {_GEN_143,_GEN_141,_GEN_139,_GEN_137,_GEN_135,_GEN_133,_GEN_131,_GEN_129}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_4942 = {_GEN_159,_GEN_157,_GEN_155,_GEN_153,_GEN_151,_GEN_149,_GEN_147,_GEN_145,_T_4934}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4949 = {_GEN_175,_GEN_173,_GEN_171,_GEN_169,_GEN_167,_GEN_165,_GEN_163,_GEN_161}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_4958 = {_GEN_191,_GEN_189,_GEN_187,_GEN_185,_GEN_183,_GEN_181,_GEN_179,_GEN_177,_T_4949,_T_4942}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4965 = {_GEN_207,_GEN_205,_GEN_203,_GEN_201,_GEN_199,_GEN_197,_GEN_195,_GEN_193}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_4973 = {_GEN_223,_GEN_221,_GEN_219,_GEN_217,_GEN_215,_GEN_213,_GEN_211,_GEN_209,_T_4965}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4980 = {_GEN_239,_GEN_237,_GEN_235,_GEN_233,_GEN_231,_GEN_229,_GEN_227,_GEN_225}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_4989 = {_GEN_255,_GEN_253,_GEN_251,_GEN_249,_GEN_247,_GEN_245,_GEN_243,_GEN_241,_T_4980,_T_4973}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_4998 = {_GEN_271,_GEN_269,_GEN_267,_GEN_265,_GEN_263,_GEN_261,_GEN_259,_GEN_257}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_5006 = {_GEN_287,_GEN_285,_GEN_283,_GEN_281,_GEN_279,_GEN_277,_GEN_275,_GEN_273,_T_4998}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5013 = {_GEN_303,_GEN_301,_GEN_299,_GEN_297,_GEN_295,_GEN_293,_GEN_291,_GEN_289}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_5022 = {_GEN_319,_GEN_317,_GEN_315,_GEN_313,_GEN_311,_GEN_309,_GEN_307,_GEN_305,_T_5013,_T_5006}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5029 = {_GEN_335,_GEN_333,_GEN_331,_GEN_329,_GEN_327,_GEN_325,_GEN_323,_GEN_321}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_5037 = {_GEN_351,_GEN_349,_GEN_347,_GEN_345,_GEN_343,_GEN_341,_GEN_339,_GEN_337,_T_5029}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5044 = {_GEN_367,_GEN_365,_GEN_363,_GEN_361,_GEN_359,_GEN_357,_GEN_355,_GEN_353}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_5053 = {_GEN_383,_GEN_381,_GEN_379,_GEN_377,_GEN_375,_GEN_373,_GEN_371,_GEN_369,_T_5044,_T_5037}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5061 = {_GEN_399,_GEN_397,_GEN_395,_GEN_393,_GEN_391,_GEN_389,_GEN_387,_GEN_385}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_5069 = {_GEN_415,_GEN_413,_GEN_411,_GEN_409,_GEN_407,_GEN_405,_GEN_403,_GEN_401,_T_5061}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5076 = {_GEN_431,_GEN_429,_GEN_427,_GEN_425,_GEN_423,_GEN_421,_GEN_419,_GEN_417}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_5085 = {_GEN_447,_GEN_445,_GEN_443,_GEN_441,_GEN_439,_GEN_437,_GEN_435,_GEN_433,_T_5076,_T_5069}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5092 = {_GEN_463,_GEN_461,_GEN_459,_GEN_457,_GEN_455,_GEN_453,_GEN_451,_GEN_449}; // @[ConwaylifeBetter.scala 42:19]
  wire [15:0] _T_5100 = {_GEN_479,_GEN_477,_GEN_475,_GEN_473,_GEN_471,_GEN_469,_GEN_467,_GEN_465,_T_5092}; // @[ConwaylifeBetter.scala 42:19]
  wire [7:0] _T_5107 = {_GEN_495,_GEN_493,_GEN_491,_GEN_489,_GEN_487,_GEN_485,_GEN_483,_GEN_481}; // @[ConwaylifeBetter.scala 42:19]
  wire [31:0] _T_5116 = {_GEN_511,_GEN_509,_GEN_507,_GEN_505,_GEN_503,_GEN_501,_GEN_499,_GEN_497,_T_5107,_T_5100}; // @[ConwaylifeBetter.scala 42:19]
  wire [255:0] _T_5119 = {_T_5116,_T_5085,_T_5053,_T_5022,_T_4989,_T_4958,_T_4926,_T_4895}; // @[ConwaylifeBetter.scala 42:19]
  assign io_q = regs; // @[ConwaylifeBetter.scala 44:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  regs = _RAND_0[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_load) begin
      regs <= io_data;
    end else begin
      regs <= _T_5119;
    end
  end
endmodule
