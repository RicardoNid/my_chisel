module CORDIC_tb;

  reg           clock;
  reg           reset;
  reg  [19 : 0] io_dataInX;
  reg  [19 : 0] io_dataInY;
  wire [49 : 0] io_dataOutX;
  wire [49 : 0] io_dataOutPhase;

  CORDIC dut (
    .clock(clock),
    .reset(reset),
    .io_dataInX(io_dataInX),
    .io_dataInY(io_dataInY),
    .io_dataOutX(io_dataOutX),
    .io_dataOutPhase(io_dataOutPhase)
  );

  initial begin
    clock      = 0;
    reset      = 0;
    io_dataInX = 0;
    io_dataInY = 0;

    #10;
    io_dataInX = 20'b11000000000000000000;
    io_dataInY = 20'b00000000000000000000;
    #10;
    io_dataInX = 20'b11000000000101100111;
    io_dataInY = 20'b11111100101001101000;
    #10;
    io_dataInX = 20'b11000000010110011100;
    io_dataInY = 20'b11111001010011110110;
    #10;
    io_dataInX = 20'b11000000110010011011;
    io_dataInY = 20'b11110101111111010000;
    #10;
    io_dataInX = 20'b11000001011001100000;
    io_dataInY = 20'b11110010101100011001;
    #10;
    io_dataInX = 20'b11000010001011100100;
    io_dataInY = 20'b11101111011011111000;
    #10;
    io_dataInX = 20'b11000011001000011110;
    io_dataInY = 20'b11101100001110010001;
    #10;
    io_dataInX = 20'b11000100010000000011;
    io_dataInY = 20'b11101001000100001000;
    #10;
    io_dataInX = 20'b11000101100010001000;
    io_dataInY = 20'b11100101111110000000;
    #10;
    io_dataInX = 20'b11000110111110011100;
    io_dataInY = 20'b11100010111100011101;
    #10;
    io_dataInX = 20'b11001000100100110001;
    io_dataInY = 20'b11100000000000000000;
    #10;
    io_dataInX = 20'b11001010010100110100;
    io_dataInY = 20'b11011101001001001010;
    #10;
    io_dataInX = 20'b11001100001110010001;
    io_dataInY = 20'b11011010011000011100;
    #10;
    io_dataInX = 20'b11001110010000110100;
    io_dataInY = 20'b11010111101110010011;
    #10;
    io_dataInX = 20'b11010000011100000101;
    io_dataInY = 20'b11010101001011001111;
    #10;
    io_dataInX = 20'b11010010101111101100;
    io_dataInY = 20'b11010010101111101100;
    #10;
    io_dataInX = 20'b11010101001011001111;
    io_dataInY = 20'b11010000011100000101;
    #10;
    io_dataInX = 20'b11010111101110010011;
    io_dataInY = 20'b11001110010000110100;
    #10;
    io_dataInX = 20'b11011010011000011100;
    io_dataInY = 20'b11001100001110010001;
    #10;
    io_dataInX = 20'b11011101001001001010;
    io_dataInY = 20'b11001010010100110100;
    #10;
    io_dataInX = 20'b11100000000000000000;
    io_dataInY = 20'b11001000100100110001;
    #10;
    io_dataInX = 20'b11100010111100011101;
    io_dataInY = 20'b11000110111110011100;
    #10;
    io_dataInX = 20'b11100101111110000000;
    io_dataInY = 20'b11000101100010001000;
    #10;
    io_dataInX = 20'b11101001000100001000;
    io_dataInY = 20'b11000100010000000011;
    #10;
    io_dataInX = 20'b11101100001110010001;
    io_dataInY = 20'b11000011001000011110;
    #10;
    io_dataInX = 20'b11101111011011111000;
    io_dataInY = 20'b11000010001011100100;
    #10;
    io_dataInX = 20'b11110010101100011001;
    io_dataInY = 20'b11000001011001100000;
    #10;
    io_dataInX = 20'b11110101111111010000;
    io_dataInY = 20'b11000000110010011011;
    #10;
    io_dataInX = 20'b11111001010011110110;
    io_dataInY = 20'b11000000010110011100;
    #10;
    io_dataInX = 20'b11111100101001101000;
    io_dataInY = 20'b11000000000101100111;
    #10;
    io_dataInX = 20'b00000000000000000000;
    io_dataInY = 20'b11000000000000000000;
    #10;
    io_dataInX = 20'b00000011010110011000;
    io_dataInY = 20'b11000000000101100111;
    #10;
    io_dataInX = 20'b00000110101100001010;
    io_dataInY = 20'b11000000010110011100;
    #10;
    io_dataInX = 20'b00001010000000110000;
    io_dataInY = 20'b11000000110010011011;
    #10;
    io_dataInX = 20'b00001101010011100111;
    io_dataInY = 20'b11000001011001100000;
    #10;
    io_dataInX = 20'b00010000100100001000;
    io_dataInY = 20'b11000010001011100100;
    #10;
    io_dataInX = 20'b00010011110001101111;
    io_dataInY = 20'b11000011001000011110;
    #10;
    io_dataInX = 20'b00010110111011111000;
    io_dataInY = 20'b11000100010000000011;
    #10;
    io_dataInX = 20'b00011010000010000000;
    io_dataInY = 20'b11000101100010001000;
    #10;
    io_dataInX = 20'b00011101000011100011;
    io_dataInY = 20'b11000110111110011100;
    #10;
    io_dataInX = 20'b00100000000000000000;
    io_dataInY = 20'b11001000100100110001;
    #10;
    io_dataInX = 20'b00100010110110110110;
    io_dataInY = 20'b11001010010100110100;
    #10;
    io_dataInX = 20'b00100101100111100100;
    io_dataInY = 20'b11001100001110010001;
    #10;
    io_dataInX = 20'b00101000010001101101;
    io_dataInY = 20'b11001110010000110100;
    #10;
    io_dataInX = 20'b00101010110100110001;
    io_dataInY = 20'b11010000011100000101;
    #10;
    io_dataInX = 20'b00101101010000010100;
    io_dataInY = 20'b11010010101111101100;
    #10;
    io_dataInX = 20'b00101111100011111011;
    io_dataInY = 20'b11010101001011001111;
    #10;
    io_dataInX = 20'b00110001101111001100;
    io_dataInY = 20'b11010111101110010011;
    #10;
    io_dataInX = 20'b00110011110001101111;
    io_dataInY = 20'b11011010011000011100;
    #10;
    io_dataInX = 20'b00110101101011001100;
    io_dataInY = 20'b11011101001001001010;
    #10;
    io_dataInX = 20'b00110111011011001111;
    io_dataInY = 20'b11100000000000000000;
    #10;
    io_dataInX = 20'b00111001000001100100;
    io_dataInY = 20'b11100010111100011101;
    #10;
    io_dataInX = 20'b00111010011101111000;
    io_dataInY = 20'b11100101111110000000;
    #10;
    io_dataInX = 20'b00111011101111111101;
    io_dataInY = 20'b11101001000100001000;
    #10;
    io_dataInX = 20'b00111100110111100010;
    io_dataInY = 20'b11101100001110010001;
    #10;
    io_dataInX = 20'b00111101110100011100;
    io_dataInY = 20'b11101111011011111000;
    #10;
    io_dataInX = 20'b00111110100110100000;
    io_dataInY = 20'b11110010101100011001;
    #10;
    io_dataInX = 20'b00111111001101100101;
    io_dataInY = 20'b11110101111111010000;
    #10;
    io_dataInX = 20'b00111111101001100100;
    io_dataInY = 20'b11111001010011110110;
    #10;
    io_dataInX = 20'b00111111111010011001;
    io_dataInY = 20'b11111100101001101000;
    #10;
    io_dataInX = 20'b01000000000000000000;
    io_dataInY = 20'b00000000000000000000;
    #10;
    io_dataInX = 20'b00111111111010011001;
    io_dataInY = 20'b00000011010110011000;
    #10;
    io_dataInX = 20'b00111111101001100100;
    io_dataInY = 20'b00000110101100001010;
    #10;
    io_dataInX = 20'b00111111001101100101;
    io_dataInY = 20'b00001010000000110000;
    #10;
    io_dataInX = 20'b00111110100110100000;
    io_dataInY = 20'b00001101010011100111;
    #10;
    io_dataInX = 20'b00111101110100011100;
    io_dataInY = 20'b00010000100100001000;
    #10;
    io_dataInX = 20'b00111100110111100010;
    io_dataInY = 20'b00010011110001101111;
    #10;
    io_dataInX = 20'b00111011101111111101;
    io_dataInY = 20'b00010110111011111000;
    #10;
    io_dataInX = 20'b00111010011101111000;
    io_dataInY = 20'b00011010000010000000;
    #10;
    io_dataInX = 20'b00111001000001100100;
    io_dataInY = 20'b00011101000011100011;
    #10;
    io_dataInX = 20'b00110111011011001111;
    io_dataInY = 20'b00100000000000000000;
    #10;
    io_dataInX = 20'b00110101101011001100;
    io_dataInY = 20'b00100010110110110110;
    #10;
    io_dataInX = 20'b00110011110001101111;
    io_dataInY = 20'b00100101100111100100;
    #10;
    io_dataInX = 20'b00110001101111001100;
    io_dataInY = 20'b00101000010001101101;
    #10;
    io_dataInX = 20'b00101111100011111011;
    io_dataInY = 20'b00101010110100110001;
    #10;
    io_dataInX = 20'b00101101010000010100;
    io_dataInY = 20'b00101101010000010100;
    #10;
    io_dataInX = 20'b00101010110100110001;
    io_dataInY = 20'b00101111100011111011;
    #10;
    io_dataInX = 20'b00101000010001101101;
    io_dataInY = 20'b00110001101111001100;
    #10;
    io_dataInX = 20'b00100101100111100100;
    io_dataInY = 20'b00110011110001101111;
    #10;
    io_dataInX = 20'b00100010110110110110;
    io_dataInY = 20'b00110101101011001100;
    #10;
    io_dataInX = 20'b00100000000000000000;
    io_dataInY = 20'b00110111011011001111;
    #10;
    io_dataInX = 20'b00011101000011100011;
    io_dataInY = 20'b00111001000001100100;
    #10;
    io_dataInX = 20'b00011010000010000000;
    io_dataInY = 20'b00111010011101111000;
    #10;
    io_dataInX = 20'b00010110111011111000;
    io_dataInY = 20'b00111011101111111101;
    #10;
    io_dataInX = 20'b00010011110001101111;
    io_dataInY = 20'b00111100110111100010;
    #10;
    io_dataInX = 20'b00010000100100001000;
    io_dataInY = 20'b00111101110100011100;
    #10;
    io_dataInX = 20'b00001101010011100111;
    io_dataInY = 20'b00111110100110100000;
    #10;
    io_dataInX = 20'b00001010000000110000;
    io_dataInY = 20'b00111111001101100101;
    #10;
    io_dataInX = 20'b00000110101100001010;
    io_dataInY = 20'b00111111101001100100;
    #10;
    io_dataInX = 20'b00000011010110011000;
    io_dataInY = 20'b00111111111010011001;
    #10;
    io_dataInX = 20'b00000000000000000000;
    io_dataInY = 20'b01000000000000000000;
    #10;
    io_dataInX = 20'b11111100101001101000;
    io_dataInY = 20'b00111111111010011001;
    #10;
    io_dataInX = 20'b11111001010011110110;
    io_dataInY = 20'b00111111101001100100;
    #10;
    io_dataInX = 20'b11110101111111010000;
    io_dataInY = 20'b00111111001101100101;
    #10;
    io_dataInX = 20'b11110010101100011001;
    io_dataInY = 20'b00111110100110100000;
    #10;
    io_dataInX = 20'b11101111011011111000;
    io_dataInY = 20'b00111101110100011100;
    #10;
    io_dataInX = 20'b11101100001110010001;
    io_dataInY = 20'b00111100110111100010;
    #10;
    io_dataInX = 20'b11101001000100001000;
    io_dataInY = 20'b00111011101111111101;
    #10;
    io_dataInX = 20'b11100101111110000000;
    io_dataInY = 20'b00111010011101111000;
    #10;
    io_dataInX = 20'b11100010111100011101;
    io_dataInY = 20'b00111001000001100100;
    #10;
    io_dataInX = 20'b11100000000000000000;
    io_dataInY = 20'b00110111011011001111;
    #10;
    io_dataInX = 20'b11011101001001001010;
    io_dataInY = 20'b00110101101011001100;
    #10;
    io_dataInX = 20'b11011010011000011100;
    io_dataInY = 20'b00110011110001101111;
    #10;
    io_dataInX = 20'b11010111101110010011;
    io_dataInY = 20'b00110001101111001100;
    #10;
    io_dataInX = 20'b11010101001011001111;
    io_dataInY = 20'b00101111100011111011;
    #10;
    io_dataInX = 20'b11010010101111101100;
    io_dataInY = 20'b00101101010000010100;
    #10;
    io_dataInX = 20'b11010000011100000101;
    io_dataInY = 20'b00101010110100110001;
    #10;
    io_dataInX = 20'b11001110010000110100;
    io_dataInY = 20'b00101000010001101101;
    #10;
    io_dataInX = 20'b11001100001110010001;
    io_dataInY = 20'b00100101100111100100;
    #10;
    io_dataInX = 20'b11001010010100110100;
    io_dataInY = 20'b00100010110110110110;
    #10;
    io_dataInX = 20'b11001000100100110001;
    io_dataInY = 20'b00100000000000000000;
    #10;
    io_dataInX = 20'b11000110111110011100;
    io_dataInY = 20'b00011101000011100011;
    #10;
    io_dataInX = 20'b11000101100010001000;
    io_dataInY = 20'b00011010000010000000;
    #10;
    io_dataInX = 20'b11000100010000000011;
    io_dataInY = 20'b00010110111011111000;
    #10;
    io_dataInX = 20'b11000011001000011110;
    io_dataInY = 20'b00010011110001101111;
    #10;
    io_dataInX = 20'b11000010001011100100;
    io_dataInY = 20'b00010000100100001000;
    #10;
    io_dataInX = 20'b11000001011001100000;
    io_dataInY = 20'b00001101010011100111;
    #10;
    io_dataInX = 20'b11000000110010011011;
    io_dataInY = 20'b00001010000000110000;
    #10;
    io_dataInX = 20'b11000000010110011100;
    io_dataInY = 20'b00000110101100001010;
    #10;
    io_dataInX = 20'b11000000000101100111;
    io_dataInY = 20'b00000011010110011000;

    #10;
    io_dataInX = 20'b10100000000000000000;
    io_dataInY = 20'b00000000000000000000;
    #10;
    io_dataInX = 20'b10100000001000011011;
    io_dataInY = 20'b00000101000001100011;
    #10;
    io_dataInX = 20'b10100000100001101010;
    io_dataInY = 20'b00001010000010001110;
    #10;
    io_dataInX = 20'b10100001001011101001;
    io_dataInY = 20'b00001111000001001001;
    #10;
    io_dataInX = 20'b10100010000110010001;
    io_dataInY = 20'b00010011111101011010;
    #10;
    io_dataInX = 20'b10100011010001010111;
    io_dataInY = 20'b00011000110110001100;
    #10;
    io_dataInX = 20'b10100100101100101101;
    io_dataInY = 20'b00011101101010100110;
    #10;
    io_dataInX = 20'b10100110011000000101;
    io_dataInY = 20'b00100010011001110100;
    #10;
    io_dataInX = 20'b10101000010011001011;
    io_dataInY = 20'b00100111000010111111;
    #10;
    io_dataInX = 20'b10101010011101101010;
    io_dataInY = 20'b00101011100101010100;
    #10;
    io_dataInX = 20'b10101100110111001001;
    io_dataInY = 20'b00110000000000000000;
    #10;
    io_dataInX = 20'b10101111011111001101;
    io_dataInY = 20'b00110100010010010001;
    #10;
    io_dataInX = 20'b10110010010101011010;
    io_dataInY = 20'b00111000011011010111;
    #10;
    io_dataInX = 20'b10110101011001001110;
    io_dataInY = 20'b00111100011010100011;
    #10;
    io_dataInX = 20'b10111000101010001000;
    io_dataInY = 20'b01000000001111001001;
    #10;
    io_dataInX = 20'b10111100000111100010;
    io_dataInY = 20'b01000011111000011110;
    #10;
    io_dataInX = 20'b10111111110000110111;
    io_dataInY = 20'b01000111010101111000;
    #10;
    io_dataInX = 20'b11000011100101011101;
    io_dataInY = 20'b01001010100110110010;
    #10;
    io_dataInX = 20'b11000111100100101001;
    io_dataInY = 20'b01001101101010100110;
    #10;
    io_dataInX = 20'b11001011101101101111;
    io_dataInY = 20'b01010000100000110011;
    #10;
    io_dataInX = 20'b11010000000000000000;
    io_dataInY = 20'b01010011001000110111;
    #10;
    io_dataInX = 20'b11010100011010101100;
    io_dataInY = 20'b01010101100010010110;
    #10;
    io_dataInX = 20'b11011000111101000001;
    io_dataInY = 20'b01010111101100110101;
    #10;
    io_dataInX = 20'b11011101100110001100;
    io_dataInY = 20'b01011001100111111011;
    #10;
    io_dataInX = 20'b11100010010101011010;
    io_dataInY = 20'b01011011010011010011;
    #10;
    io_dataInX = 20'b11100111001001110100;
    io_dataInY = 20'b01011100101110101001;
    #10;
    io_dataInX = 20'b11101100000010100110;
    io_dataInY = 20'b01011101111001101111;
    #10;
    io_dataInX = 20'b11110000111110110111;
    io_dataInY = 20'b01011110110100010111;
    #10;
    io_dataInX = 20'b11110101111101110010;
    io_dataInY = 20'b01011111011110010110;
    #10;
    io_dataInX = 20'b11111010111110011101;
    io_dataInY = 20'b01011111110111100101;
    #10;
    io_dataInX = 20'b00000000000000000000;
    io_dataInY = 20'b01100000000000000000;
    #10;
    io_dataInX = 20'b00000101000001100011;
    io_dataInY = 20'b01011111110111100101;
    #10;
    io_dataInX = 20'b00001010000010001110;
    io_dataInY = 20'b01011111011110010110;
    #10;
    io_dataInX = 20'b00001111000001001001;
    io_dataInY = 20'b01011110110100010111;
    #10;
    io_dataInX = 20'b00010011111101011010;
    io_dataInY = 20'b01011101111001101111;
    #10;
    io_dataInX = 20'b00011000110110001100;
    io_dataInY = 20'b01011100101110101001;
    #10;
    io_dataInX = 20'b00011101101010100110;
    io_dataInY = 20'b01011011010011010011;
    #10;
    io_dataInX = 20'b00100010011001110100;
    io_dataInY = 20'b01011001100111111011;
    #10;
    io_dataInX = 20'b00100111000010111111;
    io_dataInY = 20'b01010111101100110101;
    #10;
    io_dataInX = 20'b00101011100101010100;
    io_dataInY = 20'b01010101100010010110;
    #10;
    io_dataInX = 20'b00110000000000000000;
    io_dataInY = 20'b01010011001000110111;
    #10;
    io_dataInX = 20'b00110100010010010001;
    io_dataInY = 20'b01010000100000110011;
    #10;
    io_dataInX = 20'b00111000011011010111;
    io_dataInY = 20'b01001101101010100110;
    #10;
    io_dataInX = 20'b00111100011010100011;
    io_dataInY = 20'b01001010100110110010;
    #10;
    io_dataInX = 20'b01000000001111001001;
    io_dataInY = 20'b01000111010101111000;
    #10;
    io_dataInX = 20'b01000011111000011110;
    io_dataInY = 20'b01000011111000011110;
    #10;
    io_dataInX = 20'b01000111010101111000;
    io_dataInY = 20'b01000000001111001001;
    #10;
    io_dataInX = 20'b01001010100110110010;
    io_dataInY = 20'b00111100011010100011;
    #10;
    io_dataInX = 20'b01001101101010100110;
    io_dataInY = 20'b00111000011011010111;
    #10;
    io_dataInX = 20'b01010000100000110011;
    io_dataInY = 20'b00110100010010010001;
    #10;
    io_dataInX = 20'b01010011001000110111;
    io_dataInY = 20'b00110000000000000000;
    #10;
    io_dataInX = 20'b01010101100010010110;
    io_dataInY = 20'b00101011100101010100;
    #10;
    io_dataInX = 20'b01010111101100110101;
    io_dataInY = 20'b00100111000010111111;
    #10;
    io_dataInX = 20'b01011001100111111011;
    io_dataInY = 20'b00100010011001110100;
    #10;
    io_dataInX = 20'b01011011010011010011;
    io_dataInY = 20'b00011101101010100110;
    #10;
    io_dataInX = 20'b01011100101110101001;
    io_dataInY = 20'b00011000110110001100;
    #10;
    io_dataInX = 20'b01011101111001101111;
    io_dataInY = 20'b00010011111101011010;
    #10;
    io_dataInX = 20'b01011110110100010111;
    io_dataInY = 20'b00001111000001001001;
    #10;
    io_dataInX = 20'b01011111011110010110;
    io_dataInY = 20'b00001010000010001110;
    #10;
    io_dataInX = 20'b01011111110111100101;
    io_dataInY = 20'b00000101000001100011;
    #10;
    io_dataInX = 20'b01100000000000000000;
    io_dataInY = 20'b00000000000000000000;
    #10;
    io_dataInX = 20'b01011111110111100101;
    io_dataInY = 20'b11111010111110011101;
    #10;
    io_dataInX = 20'b01011111011110010110;
    io_dataInY = 20'b11110101111101110010;
    #10;
    io_dataInX = 20'b01011110110100010111;
    io_dataInY = 20'b11110000111110110111;
    #10;
    io_dataInX = 20'b01011101111001101111;
    io_dataInY = 20'b11101100000010100110;
    #10;
    io_dataInX = 20'b01011100101110101001;
    io_dataInY = 20'b11100111001001110100;
    #10;
    io_dataInX = 20'b01011011010011010011;
    io_dataInY = 20'b11100010010101011010;
    #10;
    io_dataInX = 20'b01011001100111111011;
    io_dataInY = 20'b11011101100110001100;
    #10;
    io_dataInX = 20'b01010111101100110101;
    io_dataInY = 20'b11011000111101000001;
    #10;
    io_dataInX = 20'b01010101100010010110;
    io_dataInY = 20'b11010100011010101100;
    #10;
    io_dataInX = 20'b01010011001000110111;
    io_dataInY = 20'b11010000000000000000;
    #10;
    io_dataInX = 20'b01010000100000110011;
    io_dataInY = 20'b11001011101101101111;
    #10;
    io_dataInX = 20'b01001101101010100110;
    io_dataInY = 20'b11000111100100101001;
    #10;
    io_dataInX = 20'b01001010100110110010;
    io_dataInY = 20'b11000011100101011101;
    #10;
    io_dataInX = 20'b01000111010101111000;
    io_dataInY = 20'b10111111110000110111;
    #10;
    io_dataInX = 20'b01000011111000011110;
    io_dataInY = 20'b10111100000111100010;
    #10;
    io_dataInX = 20'b01000000001111001001;
    io_dataInY = 20'b10111000101010001000;
    #10;
    io_dataInX = 20'b00111100011010100011;
    io_dataInY = 20'b10110101011001001110;
    #10;
    io_dataInX = 20'b00111000011011010111;
    io_dataInY = 20'b10110010010101011010;
    #10;
    io_dataInX = 20'b00110100010010010001;
    io_dataInY = 20'b10101111011111001101;
    #10;
    io_dataInX = 20'b00110000000000000000;
    io_dataInY = 20'b10101100110111001001;
    #10;
    io_dataInX = 20'b00101011100101010100;
    io_dataInY = 20'b10101010011101101010;
    #10;
    io_dataInX = 20'b00100111000010111111;
    io_dataInY = 20'b10101000010011001011;
    #10;
    io_dataInX = 20'b00100010011001110100;
    io_dataInY = 20'b10100110011000000101;
    #10;
    io_dataInX = 20'b00011101101010100110;
    io_dataInY = 20'b10100100101100101101;
    #10;
    io_dataInX = 20'b00011000110110001100;
    io_dataInY = 20'b10100011010001010111;
    #10;
    io_dataInX = 20'b00010011111101011010;
    io_dataInY = 20'b10100010000110010001;
    #10;
    io_dataInX = 20'b00001111000001001001;
    io_dataInY = 20'b10100001001011101001;
    #10;
    io_dataInX = 20'b00001010000010001110;
    io_dataInY = 20'b10100000100001101010;
    #10;
    io_dataInX = 20'b00000101000001100011;
    io_dataInY = 20'b10100000001000011011;
    #10;
    io_dataInX = 20'b00000000000000000000;
    io_dataInY = 20'b10100000000000000000;
    #10;
    io_dataInX = 20'b11111010111110011101;
    io_dataInY = 20'b10100000001000011011;
    #10;
    io_dataInX = 20'b11110101111101110010;
    io_dataInY = 20'b10100000100001101010;
    #10;
    io_dataInX = 20'b11110000111110110111;
    io_dataInY = 20'b10100001001011101001;
    #10;
    io_dataInX = 20'b11101100000010100110;
    io_dataInY = 20'b10100010000110010001;
    #10;
    io_dataInX = 20'b11100111001001110100;
    io_dataInY = 20'b10100011010001010111;
    #10;
    io_dataInX = 20'b11100010010101011010;
    io_dataInY = 20'b10100100101100101101;
    #10;
    io_dataInX = 20'b11011101100110001100;
    io_dataInY = 20'b10100110011000000101;
    #10;
    io_dataInX = 20'b11011000111101000001;
    io_dataInY = 20'b10101000010011001011;
    #10;
    io_dataInX = 20'b11010100011010101100;
    io_dataInY = 20'b10101010011101101010;
    #10;
    io_dataInX = 20'b11010000000000000000;
    io_dataInY = 20'b10101100110111001001;
    #10;
    io_dataInX = 20'b11001011101101101111;
    io_dataInY = 20'b10101111011111001101;
    #10;
    io_dataInX = 20'b11000111100100101001;
    io_dataInY = 20'b10110010010101011010;
    #10;
    io_dataInX = 20'b11000011100101011101;
    io_dataInY = 20'b10110101011001001110;
    #10;
    io_dataInX = 20'b10111111110000110111;
    io_dataInY = 20'b10111000101010001000;
    #10;
    io_dataInX = 20'b10111100000111100010;
    io_dataInY = 20'b10111100000111100010;
    #10;
    io_dataInX = 20'b10111000101010001000;
    io_dataInY = 20'b10111111110000110111;
    #10;
    io_dataInX = 20'b10110101011001001110;
    io_dataInY = 20'b11000011100101011101;
    #10;
    io_dataInX = 20'b10110010010101011010;
    io_dataInY = 20'b11000111100100101001;
    #10;
    io_dataInX = 20'b10101111011111001101;
    io_dataInY = 20'b11001011101101101111;
    #10;
    io_dataInX = 20'b10101100110111001001;
    io_dataInY = 20'b11010000000000000000;
    #10;
    io_dataInX = 20'b10101010011101101010;
    io_dataInY = 20'b11010100011010101100;
    #10;
    io_dataInX = 20'b10101000010011001011;
    io_dataInY = 20'b11011000111101000001;
    #10;
    io_dataInX = 20'b10100110011000000101;
    io_dataInY = 20'b11011101100110001100;
    #10;
    io_dataInX = 20'b10100100101100101101;
    io_dataInY = 20'b11100010010101011010;
    #10;
    io_dataInX = 20'b10100011010001010111;
    io_dataInY = 20'b11100111001001110100;
    #10;
    io_dataInX = 20'b10100010000110010001;
    io_dataInY = 20'b11101100000010100110;
    #10;
    io_dataInX = 20'b10100001001011101001;
    io_dataInY = 20'b11110000111110110111;
    #10;
    io_dataInX = 20'b10100000100001101010;
    io_dataInY = 20'b11110101111101110010;
    #10;
    io_dataInX = 20'b10100000001000011011;
    io_dataInY = 20'b11111010111110011101;


    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;
    #10;



  end

  always
    #5 clock = ! clock;

endmodule