module Conwaylife(
  input          clock,
  input          reset,
  input          io_load,
  input  [255:0] io_data,
  output [255:0] io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg  regs_0_0; // @[Conwaylife.scala 12:17]
  reg  regs_0_1; // @[Conwaylife.scala 12:17]
  reg  regs_0_2; // @[Conwaylife.scala 12:17]
  reg  regs_0_3; // @[Conwaylife.scala 12:17]
  reg  regs_0_4; // @[Conwaylife.scala 12:17]
  reg  regs_0_5; // @[Conwaylife.scala 12:17]
  reg  regs_0_6; // @[Conwaylife.scala 12:17]
  reg  regs_0_7; // @[Conwaylife.scala 12:17]
  reg  regs_0_8; // @[Conwaylife.scala 12:17]
  reg  regs_0_9; // @[Conwaylife.scala 12:17]
  reg  regs_0_10; // @[Conwaylife.scala 12:17]
  reg  regs_0_11; // @[Conwaylife.scala 12:17]
  reg  regs_0_12; // @[Conwaylife.scala 12:17]
  reg  regs_0_13; // @[Conwaylife.scala 12:17]
  reg  regs_0_14; // @[Conwaylife.scala 12:17]
  reg  regs_0_15; // @[Conwaylife.scala 12:17]
  reg  regs_1_0; // @[Conwaylife.scala 12:17]
  reg  regs_1_1; // @[Conwaylife.scala 12:17]
  reg  regs_1_2; // @[Conwaylife.scala 12:17]
  reg  regs_1_3; // @[Conwaylife.scala 12:17]
  reg  regs_1_4; // @[Conwaylife.scala 12:17]
  reg  regs_1_5; // @[Conwaylife.scala 12:17]
  reg  regs_1_6; // @[Conwaylife.scala 12:17]
  reg  regs_1_7; // @[Conwaylife.scala 12:17]
  reg  regs_1_8; // @[Conwaylife.scala 12:17]
  reg  regs_1_9; // @[Conwaylife.scala 12:17]
  reg  regs_1_10; // @[Conwaylife.scala 12:17]
  reg  regs_1_11; // @[Conwaylife.scala 12:17]
  reg  regs_1_12; // @[Conwaylife.scala 12:17]
  reg  regs_1_13; // @[Conwaylife.scala 12:17]
  reg  regs_1_14; // @[Conwaylife.scala 12:17]
  reg  regs_1_15; // @[Conwaylife.scala 12:17]
  reg  regs_2_0; // @[Conwaylife.scala 12:17]
  reg  regs_2_1; // @[Conwaylife.scala 12:17]
  reg  regs_2_2; // @[Conwaylife.scala 12:17]
  reg  regs_2_3; // @[Conwaylife.scala 12:17]
  reg  regs_2_4; // @[Conwaylife.scala 12:17]
  reg  regs_2_5; // @[Conwaylife.scala 12:17]
  reg  regs_2_6; // @[Conwaylife.scala 12:17]
  reg  regs_2_7; // @[Conwaylife.scala 12:17]
  reg  regs_2_8; // @[Conwaylife.scala 12:17]
  reg  regs_2_9; // @[Conwaylife.scala 12:17]
  reg  regs_2_10; // @[Conwaylife.scala 12:17]
  reg  regs_2_11; // @[Conwaylife.scala 12:17]
  reg  regs_2_12; // @[Conwaylife.scala 12:17]
  reg  regs_2_13; // @[Conwaylife.scala 12:17]
  reg  regs_2_14; // @[Conwaylife.scala 12:17]
  reg  regs_2_15; // @[Conwaylife.scala 12:17]
  reg  regs_3_0; // @[Conwaylife.scala 12:17]
  reg  regs_3_1; // @[Conwaylife.scala 12:17]
  reg  regs_3_2; // @[Conwaylife.scala 12:17]
  reg  regs_3_3; // @[Conwaylife.scala 12:17]
  reg  regs_3_4; // @[Conwaylife.scala 12:17]
  reg  regs_3_5; // @[Conwaylife.scala 12:17]
  reg  regs_3_6; // @[Conwaylife.scala 12:17]
  reg  regs_3_7; // @[Conwaylife.scala 12:17]
  reg  regs_3_8; // @[Conwaylife.scala 12:17]
  reg  regs_3_9; // @[Conwaylife.scala 12:17]
  reg  regs_3_10; // @[Conwaylife.scala 12:17]
  reg  regs_3_11; // @[Conwaylife.scala 12:17]
  reg  regs_3_12; // @[Conwaylife.scala 12:17]
  reg  regs_3_13; // @[Conwaylife.scala 12:17]
  reg  regs_3_14; // @[Conwaylife.scala 12:17]
  reg  regs_3_15; // @[Conwaylife.scala 12:17]
  reg  regs_4_0; // @[Conwaylife.scala 12:17]
  reg  regs_4_1; // @[Conwaylife.scala 12:17]
  reg  regs_4_2; // @[Conwaylife.scala 12:17]
  reg  regs_4_3; // @[Conwaylife.scala 12:17]
  reg  regs_4_4; // @[Conwaylife.scala 12:17]
  reg  regs_4_5; // @[Conwaylife.scala 12:17]
  reg  regs_4_6; // @[Conwaylife.scala 12:17]
  reg  regs_4_7; // @[Conwaylife.scala 12:17]
  reg  regs_4_8; // @[Conwaylife.scala 12:17]
  reg  regs_4_9; // @[Conwaylife.scala 12:17]
  reg  regs_4_10; // @[Conwaylife.scala 12:17]
  reg  regs_4_11; // @[Conwaylife.scala 12:17]
  reg  regs_4_12; // @[Conwaylife.scala 12:17]
  reg  regs_4_13; // @[Conwaylife.scala 12:17]
  reg  regs_4_14; // @[Conwaylife.scala 12:17]
  reg  regs_4_15; // @[Conwaylife.scala 12:17]
  reg  regs_5_0; // @[Conwaylife.scala 12:17]
  reg  regs_5_1; // @[Conwaylife.scala 12:17]
  reg  regs_5_2; // @[Conwaylife.scala 12:17]
  reg  regs_5_3; // @[Conwaylife.scala 12:17]
  reg  regs_5_4; // @[Conwaylife.scala 12:17]
  reg  regs_5_5; // @[Conwaylife.scala 12:17]
  reg  regs_5_6; // @[Conwaylife.scala 12:17]
  reg  regs_5_7; // @[Conwaylife.scala 12:17]
  reg  regs_5_8; // @[Conwaylife.scala 12:17]
  reg  regs_5_9; // @[Conwaylife.scala 12:17]
  reg  regs_5_10; // @[Conwaylife.scala 12:17]
  reg  regs_5_11; // @[Conwaylife.scala 12:17]
  reg  regs_5_12; // @[Conwaylife.scala 12:17]
  reg  regs_5_13; // @[Conwaylife.scala 12:17]
  reg  regs_5_14; // @[Conwaylife.scala 12:17]
  reg  regs_5_15; // @[Conwaylife.scala 12:17]
  reg  regs_6_0; // @[Conwaylife.scala 12:17]
  reg  regs_6_1; // @[Conwaylife.scala 12:17]
  reg  regs_6_2; // @[Conwaylife.scala 12:17]
  reg  regs_6_3; // @[Conwaylife.scala 12:17]
  reg  regs_6_4; // @[Conwaylife.scala 12:17]
  reg  regs_6_5; // @[Conwaylife.scala 12:17]
  reg  regs_6_6; // @[Conwaylife.scala 12:17]
  reg  regs_6_7; // @[Conwaylife.scala 12:17]
  reg  regs_6_8; // @[Conwaylife.scala 12:17]
  reg  regs_6_9; // @[Conwaylife.scala 12:17]
  reg  regs_6_10; // @[Conwaylife.scala 12:17]
  reg  regs_6_11; // @[Conwaylife.scala 12:17]
  reg  regs_6_12; // @[Conwaylife.scala 12:17]
  reg  regs_6_13; // @[Conwaylife.scala 12:17]
  reg  regs_6_14; // @[Conwaylife.scala 12:17]
  reg  regs_6_15; // @[Conwaylife.scala 12:17]
  reg  regs_7_0; // @[Conwaylife.scala 12:17]
  reg  regs_7_1; // @[Conwaylife.scala 12:17]
  reg  regs_7_2; // @[Conwaylife.scala 12:17]
  reg  regs_7_3; // @[Conwaylife.scala 12:17]
  reg  regs_7_4; // @[Conwaylife.scala 12:17]
  reg  regs_7_5; // @[Conwaylife.scala 12:17]
  reg  regs_7_6; // @[Conwaylife.scala 12:17]
  reg  regs_7_7; // @[Conwaylife.scala 12:17]
  reg  regs_7_8; // @[Conwaylife.scala 12:17]
  reg  regs_7_9; // @[Conwaylife.scala 12:17]
  reg  regs_7_10; // @[Conwaylife.scala 12:17]
  reg  regs_7_11; // @[Conwaylife.scala 12:17]
  reg  regs_7_12; // @[Conwaylife.scala 12:17]
  reg  regs_7_13; // @[Conwaylife.scala 12:17]
  reg  regs_7_14; // @[Conwaylife.scala 12:17]
  reg  regs_7_15; // @[Conwaylife.scala 12:17]
  reg  regs_8_0; // @[Conwaylife.scala 12:17]
  reg  regs_8_1; // @[Conwaylife.scala 12:17]
  reg  regs_8_2; // @[Conwaylife.scala 12:17]
  reg  regs_8_3; // @[Conwaylife.scala 12:17]
  reg  regs_8_4; // @[Conwaylife.scala 12:17]
  reg  regs_8_5; // @[Conwaylife.scala 12:17]
  reg  regs_8_6; // @[Conwaylife.scala 12:17]
  reg  regs_8_7; // @[Conwaylife.scala 12:17]
  reg  regs_8_8; // @[Conwaylife.scala 12:17]
  reg  regs_8_9; // @[Conwaylife.scala 12:17]
  reg  regs_8_10; // @[Conwaylife.scala 12:17]
  reg  regs_8_11; // @[Conwaylife.scala 12:17]
  reg  regs_8_12; // @[Conwaylife.scala 12:17]
  reg  regs_8_13; // @[Conwaylife.scala 12:17]
  reg  regs_8_14; // @[Conwaylife.scala 12:17]
  reg  regs_8_15; // @[Conwaylife.scala 12:17]
  reg  regs_9_0; // @[Conwaylife.scala 12:17]
  reg  regs_9_1; // @[Conwaylife.scala 12:17]
  reg  regs_9_2; // @[Conwaylife.scala 12:17]
  reg  regs_9_3; // @[Conwaylife.scala 12:17]
  reg  regs_9_4; // @[Conwaylife.scala 12:17]
  reg  regs_9_5; // @[Conwaylife.scala 12:17]
  reg  regs_9_6; // @[Conwaylife.scala 12:17]
  reg  regs_9_7; // @[Conwaylife.scala 12:17]
  reg  regs_9_8; // @[Conwaylife.scala 12:17]
  reg  regs_9_9; // @[Conwaylife.scala 12:17]
  reg  regs_9_10; // @[Conwaylife.scala 12:17]
  reg  regs_9_11; // @[Conwaylife.scala 12:17]
  reg  regs_9_12; // @[Conwaylife.scala 12:17]
  reg  regs_9_13; // @[Conwaylife.scala 12:17]
  reg  regs_9_14; // @[Conwaylife.scala 12:17]
  reg  regs_9_15; // @[Conwaylife.scala 12:17]
  reg  regs_10_0; // @[Conwaylife.scala 12:17]
  reg  regs_10_1; // @[Conwaylife.scala 12:17]
  reg  regs_10_2; // @[Conwaylife.scala 12:17]
  reg  regs_10_3; // @[Conwaylife.scala 12:17]
  reg  regs_10_4; // @[Conwaylife.scala 12:17]
  reg  regs_10_5; // @[Conwaylife.scala 12:17]
  reg  regs_10_6; // @[Conwaylife.scala 12:17]
  reg  regs_10_7; // @[Conwaylife.scala 12:17]
  reg  regs_10_8; // @[Conwaylife.scala 12:17]
  reg  regs_10_9; // @[Conwaylife.scala 12:17]
  reg  regs_10_10; // @[Conwaylife.scala 12:17]
  reg  regs_10_11; // @[Conwaylife.scala 12:17]
  reg  regs_10_12; // @[Conwaylife.scala 12:17]
  reg  regs_10_13; // @[Conwaylife.scala 12:17]
  reg  regs_10_14; // @[Conwaylife.scala 12:17]
  reg  regs_10_15; // @[Conwaylife.scala 12:17]
  reg  regs_11_0; // @[Conwaylife.scala 12:17]
  reg  regs_11_1; // @[Conwaylife.scala 12:17]
  reg  regs_11_2; // @[Conwaylife.scala 12:17]
  reg  regs_11_3; // @[Conwaylife.scala 12:17]
  reg  regs_11_4; // @[Conwaylife.scala 12:17]
  reg  regs_11_5; // @[Conwaylife.scala 12:17]
  reg  regs_11_6; // @[Conwaylife.scala 12:17]
  reg  regs_11_7; // @[Conwaylife.scala 12:17]
  reg  regs_11_8; // @[Conwaylife.scala 12:17]
  reg  regs_11_9; // @[Conwaylife.scala 12:17]
  reg  regs_11_10; // @[Conwaylife.scala 12:17]
  reg  regs_11_11; // @[Conwaylife.scala 12:17]
  reg  regs_11_12; // @[Conwaylife.scala 12:17]
  reg  regs_11_13; // @[Conwaylife.scala 12:17]
  reg  regs_11_14; // @[Conwaylife.scala 12:17]
  reg  regs_11_15; // @[Conwaylife.scala 12:17]
  reg  regs_12_0; // @[Conwaylife.scala 12:17]
  reg  regs_12_1; // @[Conwaylife.scala 12:17]
  reg  regs_12_2; // @[Conwaylife.scala 12:17]
  reg  regs_12_3; // @[Conwaylife.scala 12:17]
  reg  regs_12_4; // @[Conwaylife.scala 12:17]
  reg  regs_12_5; // @[Conwaylife.scala 12:17]
  reg  regs_12_6; // @[Conwaylife.scala 12:17]
  reg  regs_12_7; // @[Conwaylife.scala 12:17]
  reg  regs_12_8; // @[Conwaylife.scala 12:17]
  reg  regs_12_9; // @[Conwaylife.scala 12:17]
  reg  regs_12_10; // @[Conwaylife.scala 12:17]
  reg  regs_12_11; // @[Conwaylife.scala 12:17]
  reg  regs_12_12; // @[Conwaylife.scala 12:17]
  reg  regs_12_13; // @[Conwaylife.scala 12:17]
  reg  regs_12_14; // @[Conwaylife.scala 12:17]
  reg  regs_12_15; // @[Conwaylife.scala 12:17]
  reg  regs_13_0; // @[Conwaylife.scala 12:17]
  reg  regs_13_1; // @[Conwaylife.scala 12:17]
  reg  regs_13_2; // @[Conwaylife.scala 12:17]
  reg  regs_13_3; // @[Conwaylife.scala 12:17]
  reg  regs_13_4; // @[Conwaylife.scala 12:17]
  reg  regs_13_5; // @[Conwaylife.scala 12:17]
  reg  regs_13_6; // @[Conwaylife.scala 12:17]
  reg  regs_13_7; // @[Conwaylife.scala 12:17]
  reg  regs_13_8; // @[Conwaylife.scala 12:17]
  reg  regs_13_9; // @[Conwaylife.scala 12:17]
  reg  regs_13_10; // @[Conwaylife.scala 12:17]
  reg  regs_13_11; // @[Conwaylife.scala 12:17]
  reg  regs_13_12; // @[Conwaylife.scala 12:17]
  reg  regs_13_13; // @[Conwaylife.scala 12:17]
  reg  regs_13_14; // @[Conwaylife.scala 12:17]
  reg  regs_13_15; // @[Conwaylife.scala 12:17]
  reg  regs_14_0; // @[Conwaylife.scala 12:17]
  reg  regs_14_1; // @[Conwaylife.scala 12:17]
  reg  regs_14_2; // @[Conwaylife.scala 12:17]
  reg  regs_14_3; // @[Conwaylife.scala 12:17]
  reg  regs_14_4; // @[Conwaylife.scala 12:17]
  reg  regs_14_5; // @[Conwaylife.scala 12:17]
  reg  regs_14_6; // @[Conwaylife.scala 12:17]
  reg  regs_14_7; // @[Conwaylife.scala 12:17]
  reg  regs_14_8; // @[Conwaylife.scala 12:17]
  reg  regs_14_9; // @[Conwaylife.scala 12:17]
  reg  regs_14_10; // @[Conwaylife.scala 12:17]
  reg  regs_14_11; // @[Conwaylife.scala 12:17]
  reg  regs_14_12; // @[Conwaylife.scala 12:17]
  reg  regs_14_13; // @[Conwaylife.scala 12:17]
  reg  regs_14_14; // @[Conwaylife.scala 12:17]
  reg  regs_14_15; // @[Conwaylife.scala 12:17]
  reg  regs_15_0; // @[Conwaylife.scala 12:17]
  reg  regs_15_1; // @[Conwaylife.scala 12:17]
  reg  regs_15_2; // @[Conwaylife.scala 12:17]
  reg  regs_15_3; // @[Conwaylife.scala 12:17]
  reg  regs_15_4; // @[Conwaylife.scala 12:17]
  reg  regs_15_5; // @[Conwaylife.scala 12:17]
  reg  regs_15_6; // @[Conwaylife.scala 12:17]
  reg  regs_15_7; // @[Conwaylife.scala 12:17]
  reg  regs_15_8; // @[Conwaylife.scala 12:17]
  reg  regs_15_9; // @[Conwaylife.scala 12:17]
  reg  regs_15_10; // @[Conwaylife.scala 12:17]
  reg  regs_15_11; // @[Conwaylife.scala 12:17]
  reg  regs_15_12; // @[Conwaylife.scala 12:17]
  reg  regs_15_13; // @[Conwaylife.scala 12:17]
  reg  regs_15_14; // @[Conwaylife.scala 12:17]
  reg  regs_15_15; // @[Conwaylife.scala 12:17]
  wire [1:0] _T_257 = regs_15_15 + regs_15_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1024 = {{1'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_258 = _T_257 + _GEN_1024; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1025 = {{2'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_259 = _T_258 + _GEN_1025; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1026 = {{3'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_260 = _T_259 + _GEN_1026; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1027 = {{4'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_261 = _T_260 + _GEN_1027; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1028 = {{5'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_262 = _T_261 + _GEN_1028; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1029 = {{6'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_263 = _T_262 + _GEN_1029; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1030 = {{7'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_264 = _T_263 + _GEN_1030; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1031 = {{8'd0}, regs_0_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_266 = _T_264 - _GEN_1031; // @[Conwaylife.scala 29:42]
  wire  _T_267 = _T_266 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_268 = _T_266 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_269 = _T_266 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_271 = regs_15_0 + regs_15_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1032 = {{1'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_272 = _T_271 + _GEN_1032; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1033 = {{2'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_273 = _T_272 + _GEN_1033; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1034 = {{3'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_274 = _T_273 + _GEN_1034; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1035 = {{4'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_275 = _T_274 + _GEN_1035; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1036 = {{5'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_276 = _T_275 + _GEN_1036; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1037 = {{6'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_277 = _T_276 + _GEN_1037; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1038 = {{7'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_278 = _T_277 + _GEN_1038; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1039 = {{8'd0}, regs_0_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_280 = _T_278 - _GEN_1039; // @[Conwaylife.scala 29:42]
  wire  _T_281 = _T_280 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_282 = _T_280 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_283 = _T_280 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_285 = regs_15_1 + regs_15_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1040 = {{1'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_286 = _T_285 + _GEN_1040; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1041 = {{2'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_287 = _T_286 + _GEN_1041; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1042 = {{3'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_288 = _T_287 + _GEN_1042; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1043 = {{4'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_289 = _T_288 + _GEN_1043; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1044 = {{5'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_290 = _T_289 + _GEN_1044; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1045 = {{6'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_291 = _T_290 + _GEN_1045; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1046 = {{7'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_292 = _T_291 + _GEN_1046; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1047 = {{8'd0}, regs_0_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_294 = _T_292 - _GEN_1047; // @[Conwaylife.scala 29:42]
  wire  _T_295 = _T_294 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_296 = _T_294 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_297 = _T_294 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_299 = regs_15_2 + regs_15_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1048 = {{1'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_300 = _T_299 + _GEN_1048; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1049 = {{2'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_301 = _T_300 + _GEN_1049; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1050 = {{3'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_302 = _T_301 + _GEN_1050; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1051 = {{4'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_303 = _T_302 + _GEN_1051; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1052 = {{5'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_304 = _T_303 + _GEN_1052; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1053 = {{6'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_305 = _T_304 + _GEN_1053; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1054 = {{7'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_306 = _T_305 + _GEN_1054; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1055 = {{8'd0}, regs_0_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_308 = _T_306 - _GEN_1055; // @[Conwaylife.scala 29:42]
  wire  _T_309 = _T_308 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_310 = _T_308 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_311 = _T_308 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_313 = regs_15_3 + regs_15_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1056 = {{1'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_314 = _T_313 + _GEN_1056; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1057 = {{2'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_315 = _T_314 + _GEN_1057; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1058 = {{3'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_316 = _T_315 + _GEN_1058; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1059 = {{4'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_317 = _T_316 + _GEN_1059; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1060 = {{5'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_318 = _T_317 + _GEN_1060; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1061 = {{6'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_319 = _T_318 + _GEN_1061; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1062 = {{7'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_320 = _T_319 + _GEN_1062; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1063 = {{8'd0}, regs_0_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_322 = _T_320 - _GEN_1063; // @[Conwaylife.scala 29:42]
  wire  _T_323 = _T_322 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_324 = _T_322 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_325 = _T_322 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_327 = regs_15_4 + regs_15_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1064 = {{1'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_328 = _T_327 + _GEN_1064; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1065 = {{2'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_329 = _T_328 + _GEN_1065; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1066 = {{3'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_330 = _T_329 + _GEN_1066; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1067 = {{4'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_331 = _T_330 + _GEN_1067; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1068 = {{5'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_332 = _T_331 + _GEN_1068; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1069 = {{6'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_333 = _T_332 + _GEN_1069; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1070 = {{7'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_334 = _T_333 + _GEN_1070; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1071 = {{8'd0}, regs_0_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_336 = _T_334 - _GEN_1071; // @[Conwaylife.scala 29:42]
  wire  _T_337 = _T_336 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_338 = _T_336 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_339 = _T_336 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_341 = regs_15_5 + regs_15_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1072 = {{1'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_342 = _T_341 + _GEN_1072; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1073 = {{2'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_343 = _T_342 + _GEN_1073; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1074 = {{3'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_344 = _T_343 + _GEN_1074; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1075 = {{4'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_345 = _T_344 + _GEN_1075; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1076 = {{5'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_346 = _T_345 + _GEN_1076; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1077 = {{6'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_347 = _T_346 + _GEN_1077; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1078 = {{7'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_348 = _T_347 + _GEN_1078; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1079 = {{8'd0}, regs_0_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_350 = _T_348 - _GEN_1079; // @[Conwaylife.scala 29:42]
  wire  _T_351 = _T_350 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_352 = _T_350 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_353 = _T_350 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_355 = regs_15_6 + regs_15_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1080 = {{1'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_356 = _T_355 + _GEN_1080; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1081 = {{2'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_357 = _T_356 + _GEN_1081; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1082 = {{3'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_358 = _T_357 + _GEN_1082; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1083 = {{4'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_359 = _T_358 + _GEN_1083; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1084 = {{5'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_360 = _T_359 + _GEN_1084; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1085 = {{6'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_361 = _T_360 + _GEN_1085; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1086 = {{7'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_362 = _T_361 + _GEN_1086; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1087 = {{8'd0}, regs_0_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_364 = _T_362 - _GEN_1087; // @[Conwaylife.scala 29:42]
  wire  _T_365 = _T_364 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_366 = _T_364 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_367 = _T_364 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_369 = regs_15_7 + regs_15_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1088 = {{1'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_370 = _T_369 + _GEN_1088; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1089 = {{2'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_371 = _T_370 + _GEN_1089; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1090 = {{3'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_372 = _T_371 + _GEN_1090; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1091 = {{4'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_373 = _T_372 + _GEN_1091; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1092 = {{5'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_374 = _T_373 + _GEN_1092; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1093 = {{6'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_375 = _T_374 + _GEN_1093; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1094 = {{7'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_376 = _T_375 + _GEN_1094; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1095 = {{8'd0}, regs_0_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_378 = _T_376 - _GEN_1095; // @[Conwaylife.scala 29:42]
  wire  _T_379 = _T_378 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_380 = _T_378 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_381 = _T_378 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_383 = regs_15_8 + regs_15_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1096 = {{1'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_384 = _T_383 + _GEN_1096; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1097 = {{2'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_385 = _T_384 + _GEN_1097; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1098 = {{3'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_386 = _T_385 + _GEN_1098; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1099 = {{4'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_387 = _T_386 + _GEN_1099; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1100 = {{5'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_388 = _T_387 + _GEN_1100; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1101 = {{6'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_389 = _T_388 + _GEN_1101; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1102 = {{7'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_390 = _T_389 + _GEN_1102; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1103 = {{8'd0}, regs_0_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_392 = _T_390 - _GEN_1103; // @[Conwaylife.scala 29:42]
  wire  _T_393 = _T_392 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_394 = _T_392 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_395 = _T_392 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_397 = regs_15_9 + regs_15_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1104 = {{1'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_398 = _T_397 + _GEN_1104; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1105 = {{2'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_399 = _T_398 + _GEN_1105; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1106 = {{3'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_400 = _T_399 + _GEN_1106; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1107 = {{4'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_401 = _T_400 + _GEN_1107; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1108 = {{5'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_402 = _T_401 + _GEN_1108; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1109 = {{6'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_403 = _T_402 + _GEN_1109; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1110 = {{7'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_404 = _T_403 + _GEN_1110; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1111 = {{8'd0}, regs_0_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_406 = _T_404 - _GEN_1111; // @[Conwaylife.scala 29:42]
  wire  _T_407 = _T_406 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_408 = _T_406 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_409 = _T_406 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_411 = regs_15_10 + regs_15_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1112 = {{1'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_412 = _T_411 + _GEN_1112; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1113 = {{2'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_413 = _T_412 + _GEN_1113; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1114 = {{3'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_414 = _T_413 + _GEN_1114; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1115 = {{4'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_415 = _T_414 + _GEN_1115; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1116 = {{5'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_416 = _T_415 + _GEN_1116; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1117 = {{6'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_417 = _T_416 + _GEN_1117; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1118 = {{7'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_418 = _T_417 + _GEN_1118; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1119 = {{8'd0}, regs_0_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_420 = _T_418 - _GEN_1119; // @[Conwaylife.scala 29:42]
  wire  _T_421 = _T_420 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_422 = _T_420 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_423 = _T_420 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_425 = regs_15_11 + regs_15_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1120 = {{1'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_426 = _T_425 + _GEN_1120; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1121 = {{2'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_427 = _T_426 + _GEN_1121; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1122 = {{3'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_428 = _T_427 + _GEN_1122; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1123 = {{4'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_429 = _T_428 + _GEN_1123; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1124 = {{5'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_430 = _T_429 + _GEN_1124; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1125 = {{6'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_431 = _T_430 + _GEN_1125; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1126 = {{7'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_432 = _T_431 + _GEN_1126; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1127 = {{8'd0}, regs_0_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_434 = _T_432 - _GEN_1127; // @[Conwaylife.scala 29:42]
  wire  _T_435 = _T_434 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_436 = _T_434 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_437 = _T_434 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_439 = regs_15_12 + regs_15_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1128 = {{1'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_440 = _T_439 + _GEN_1128; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1129 = {{2'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_441 = _T_440 + _GEN_1129; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1130 = {{3'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_442 = _T_441 + _GEN_1130; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1131 = {{4'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_443 = _T_442 + _GEN_1131; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1132 = {{5'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_444 = _T_443 + _GEN_1132; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1133 = {{6'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_445 = _T_444 + _GEN_1133; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1134 = {{7'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_446 = _T_445 + _GEN_1134; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1135 = {{8'd0}, regs_0_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_448 = _T_446 - _GEN_1135; // @[Conwaylife.scala 29:42]
  wire  _T_449 = _T_448 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_450 = _T_448 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_451 = _T_448 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_453 = regs_15_13 + regs_15_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1136 = {{1'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_454 = _T_453 + _GEN_1136; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1137 = {{2'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_455 = _T_454 + _GEN_1137; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1138 = {{3'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_456 = _T_455 + _GEN_1138; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1139 = {{4'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_457 = _T_456 + _GEN_1139; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1140 = {{5'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_458 = _T_457 + _GEN_1140; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1141 = {{6'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_459 = _T_458 + _GEN_1141; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1142 = {{7'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_460 = _T_459 + _GEN_1142; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1143 = {{8'd0}, regs_0_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_462 = _T_460 - _GEN_1143; // @[Conwaylife.scala 29:42]
  wire  _T_463 = _T_462 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_464 = _T_462 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_465 = _T_462 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_467 = regs_15_14 + regs_15_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1144 = {{1'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_468 = _T_467 + _GEN_1144; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1145 = {{2'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_469 = _T_468 + _GEN_1145; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1146 = {{3'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_470 = _T_469 + _GEN_1146; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1147 = {{4'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_471 = _T_470 + _GEN_1147; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1148 = {{5'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_472 = _T_471 + _GEN_1148; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1149 = {{6'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_473 = _T_472 + _GEN_1149; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1150 = {{7'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_474 = _T_473 + _GEN_1150; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1151 = {{8'd0}, regs_0_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_476 = _T_474 - _GEN_1151; // @[Conwaylife.scala 29:42]
  wire  _T_477 = _T_476 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_478 = _T_476 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_479 = _T_476 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_481 = regs_0_15 + regs_0_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1152 = {{1'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_482 = _T_481 + _GEN_1152; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1153 = {{2'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_483 = _T_482 + _GEN_1153; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1154 = {{3'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_484 = _T_483 + _GEN_1154; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1155 = {{4'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_485 = _T_484 + _GEN_1155; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1156 = {{5'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_486 = _T_485 + _GEN_1156; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1157 = {{6'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_487 = _T_486 + _GEN_1157; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1158 = {{7'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_488 = _T_487 + _GEN_1158; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1159 = {{8'd0}, regs_1_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_490 = _T_488 - _GEN_1159; // @[Conwaylife.scala 29:42]
  wire  _T_491 = _T_490 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_492 = _T_490 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_493 = _T_490 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_495 = regs_0_0 + regs_0_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1160 = {{1'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_496 = _T_495 + _GEN_1160; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1161 = {{2'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_497 = _T_496 + _GEN_1161; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1162 = {{3'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_498 = _T_497 + _GEN_1162; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1163 = {{4'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_499 = _T_498 + _GEN_1163; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1164 = {{5'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_500 = _T_499 + _GEN_1164; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1165 = {{6'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_501 = _T_500 + _GEN_1165; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1166 = {{7'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_502 = _T_501 + _GEN_1166; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1167 = {{8'd0}, regs_1_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_504 = _T_502 - _GEN_1167; // @[Conwaylife.scala 29:42]
  wire  _T_505 = _T_504 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_506 = _T_504 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_507 = _T_504 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_509 = regs_0_1 + regs_0_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1168 = {{1'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_510 = _T_509 + _GEN_1168; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1169 = {{2'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_511 = _T_510 + _GEN_1169; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1170 = {{3'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_512 = _T_511 + _GEN_1170; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1171 = {{4'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_513 = _T_512 + _GEN_1171; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1172 = {{5'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_514 = _T_513 + _GEN_1172; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1173 = {{6'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_515 = _T_514 + _GEN_1173; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1174 = {{7'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_516 = _T_515 + _GEN_1174; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1175 = {{8'd0}, regs_1_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_518 = _T_516 - _GEN_1175; // @[Conwaylife.scala 29:42]
  wire  _T_519 = _T_518 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_520 = _T_518 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_521 = _T_518 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_523 = regs_0_2 + regs_0_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1176 = {{1'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_524 = _T_523 + _GEN_1176; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1177 = {{2'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_525 = _T_524 + _GEN_1177; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1178 = {{3'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_526 = _T_525 + _GEN_1178; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1179 = {{4'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_527 = _T_526 + _GEN_1179; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1180 = {{5'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_528 = _T_527 + _GEN_1180; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1181 = {{6'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_529 = _T_528 + _GEN_1181; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1182 = {{7'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_530 = _T_529 + _GEN_1182; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1183 = {{8'd0}, regs_1_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_532 = _T_530 - _GEN_1183; // @[Conwaylife.scala 29:42]
  wire  _T_533 = _T_532 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_534 = _T_532 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_535 = _T_532 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_537 = regs_0_3 + regs_0_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1184 = {{1'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_538 = _T_537 + _GEN_1184; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1185 = {{2'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_539 = _T_538 + _GEN_1185; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1186 = {{3'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_540 = _T_539 + _GEN_1186; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1187 = {{4'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_541 = _T_540 + _GEN_1187; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1188 = {{5'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_542 = _T_541 + _GEN_1188; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1189 = {{6'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_543 = _T_542 + _GEN_1189; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1190 = {{7'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_544 = _T_543 + _GEN_1190; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1191 = {{8'd0}, regs_1_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_546 = _T_544 - _GEN_1191; // @[Conwaylife.scala 29:42]
  wire  _T_547 = _T_546 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_548 = _T_546 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_549 = _T_546 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_551 = regs_0_4 + regs_0_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1192 = {{1'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_552 = _T_551 + _GEN_1192; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1193 = {{2'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_553 = _T_552 + _GEN_1193; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1194 = {{3'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_554 = _T_553 + _GEN_1194; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1195 = {{4'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_555 = _T_554 + _GEN_1195; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1196 = {{5'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_556 = _T_555 + _GEN_1196; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1197 = {{6'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_557 = _T_556 + _GEN_1197; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1198 = {{7'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_558 = _T_557 + _GEN_1198; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1199 = {{8'd0}, regs_1_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_560 = _T_558 - _GEN_1199; // @[Conwaylife.scala 29:42]
  wire  _T_561 = _T_560 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_562 = _T_560 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_563 = _T_560 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_565 = regs_0_5 + regs_0_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1200 = {{1'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_566 = _T_565 + _GEN_1200; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1201 = {{2'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_567 = _T_566 + _GEN_1201; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1202 = {{3'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_568 = _T_567 + _GEN_1202; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1203 = {{4'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_569 = _T_568 + _GEN_1203; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1204 = {{5'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_570 = _T_569 + _GEN_1204; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1205 = {{6'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_571 = _T_570 + _GEN_1205; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1206 = {{7'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_572 = _T_571 + _GEN_1206; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1207 = {{8'd0}, regs_1_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_574 = _T_572 - _GEN_1207; // @[Conwaylife.scala 29:42]
  wire  _T_575 = _T_574 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_576 = _T_574 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_577 = _T_574 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_579 = regs_0_6 + regs_0_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1208 = {{1'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_580 = _T_579 + _GEN_1208; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1209 = {{2'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_581 = _T_580 + _GEN_1209; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1210 = {{3'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_582 = _T_581 + _GEN_1210; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1211 = {{4'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_583 = _T_582 + _GEN_1211; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1212 = {{5'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_584 = _T_583 + _GEN_1212; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1213 = {{6'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_585 = _T_584 + _GEN_1213; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1214 = {{7'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_586 = _T_585 + _GEN_1214; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1215 = {{8'd0}, regs_1_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_588 = _T_586 - _GEN_1215; // @[Conwaylife.scala 29:42]
  wire  _T_589 = _T_588 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_590 = _T_588 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_591 = _T_588 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_593 = regs_0_7 + regs_0_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1216 = {{1'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_594 = _T_593 + _GEN_1216; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1217 = {{2'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_595 = _T_594 + _GEN_1217; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1218 = {{3'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_596 = _T_595 + _GEN_1218; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1219 = {{4'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_597 = _T_596 + _GEN_1219; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1220 = {{5'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_598 = _T_597 + _GEN_1220; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1221 = {{6'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_599 = _T_598 + _GEN_1221; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1222 = {{7'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_600 = _T_599 + _GEN_1222; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1223 = {{8'd0}, regs_1_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_602 = _T_600 - _GEN_1223; // @[Conwaylife.scala 29:42]
  wire  _T_603 = _T_602 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_604 = _T_602 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_605 = _T_602 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_607 = regs_0_8 + regs_0_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1224 = {{1'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_608 = _T_607 + _GEN_1224; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1225 = {{2'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_609 = _T_608 + _GEN_1225; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1226 = {{3'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_610 = _T_609 + _GEN_1226; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1227 = {{4'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_611 = _T_610 + _GEN_1227; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1228 = {{5'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_612 = _T_611 + _GEN_1228; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1229 = {{6'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_613 = _T_612 + _GEN_1229; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1230 = {{7'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_614 = _T_613 + _GEN_1230; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1231 = {{8'd0}, regs_1_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_616 = _T_614 - _GEN_1231; // @[Conwaylife.scala 29:42]
  wire  _T_617 = _T_616 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_618 = _T_616 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_619 = _T_616 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_621 = regs_0_9 + regs_0_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1232 = {{1'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_622 = _T_621 + _GEN_1232; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1233 = {{2'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_623 = _T_622 + _GEN_1233; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1234 = {{3'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_624 = _T_623 + _GEN_1234; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1235 = {{4'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_625 = _T_624 + _GEN_1235; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1236 = {{5'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_626 = _T_625 + _GEN_1236; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1237 = {{6'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_627 = _T_626 + _GEN_1237; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1238 = {{7'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_628 = _T_627 + _GEN_1238; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1239 = {{8'd0}, regs_1_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_630 = _T_628 - _GEN_1239; // @[Conwaylife.scala 29:42]
  wire  _T_631 = _T_630 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_632 = _T_630 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_633 = _T_630 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_635 = regs_0_10 + regs_0_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1240 = {{1'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_636 = _T_635 + _GEN_1240; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1241 = {{2'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_637 = _T_636 + _GEN_1241; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1242 = {{3'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_638 = _T_637 + _GEN_1242; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1243 = {{4'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_639 = _T_638 + _GEN_1243; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1244 = {{5'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_640 = _T_639 + _GEN_1244; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1245 = {{6'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_641 = _T_640 + _GEN_1245; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1246 = {{7'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_642 = _T_641 + _GEN_1246; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1247 = {{8'd0}, regs_1_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_644 = _T_642 - _GEN_1247; // @[Conwaylife.scala 29:42]
  wire  _T_645 = _T_644 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_646 = _T_644 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_647 = _T_644 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_649 = regs_0_11 + regs_0_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1248 = {{1'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_650 = _T_649 + _GEN_1248; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1249 = {{2'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_651 = _T_650 + _GEN_1249; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1250 = {{3'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_652 = _T_651 + _GEN_1250; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1251 = {{4'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_653 = _T_652 + _GEN_1251; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1252 = {{5'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_654 = _T_653 + _GEN_1252; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1253 = {{6'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_655 = _T_654 + _GEN_1253; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1254 = {{7'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_656 = _T_655 + _GEN_1254; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1255 = {{8'd0}, regs_1_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_658 = _T_656 - _GEN_1255; // @[Conwaylife.scala 29:42]
  wire  _T_659 = _T_658 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_660 = _T_658 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_661 = _T_658 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_663 = regs_0_12 + regs_0_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1256 = {{1'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_664 = _T_663 + _GEN_1256; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1257 = {{2'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_665 = _T_664 + _GEN_1257; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1258 = {{3'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_666 = _T_665 + _GEN_1258; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1259 = {{4'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_667 = _T_666 + _GEN_1259; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1260 = {{5'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_668 = _T_667 + _GEN_1260; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1261 = {{6'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_669 = _T_668 + _GEN_1261; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1262 = {{7'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_670 = _T_669 + _GEN_1262; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1263 = {{8'd0}, regs_1_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_672 = _T_670 - _GEN_1263; // @[Conwaylife.scala 29:42]
  wire  _T_673 = _T_672 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_674 = _T_672 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_675 = _T_672 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_677 = regs_0_13 + regs_0_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1264 = {{1'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_678 = _T_677 + _GEN_1264; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1265 = {{2'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_679 = _T_678 + _GEN_1265; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1266 = {{3'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_680 = _T_679 + _GEN_1266; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1267 = {{4'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_681 = _T_680 + _GEN_1267; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1268 = {{5'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_682 = _T_681 + _GEN_1268; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1269 = {{6'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_683 = _T_682 + _GEN_1269; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1270 = {{7'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_684 = _T_683 + _GEN_1270; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1271 = {{8'd0}, regs_1_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_686 = _T_684 - _GEN_1271; // @[Conwaylife.scala 29:42]
  wire  _T_687 = _T_686 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_688 = _T_686 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_689 = _T_686 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_691 = regs_0_14 + regs_0_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1272 = {{1'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_692 = _T_691 + _GEN_1272; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1273 = {{2'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_693 = _T_692 + _GEN_1273; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1274 = {{3'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_694 = _T_693 + _GEN_1274; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1275 = {{4'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_695 = _T_694 + _GEN_1275; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1276 = {{5'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_696 = _T_695 + _GEN_1276; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1277 = {{6'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_697 = _T_696 + _GEN_1277; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1278 = {{7'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_698 = _T_697 + _GEN_1278; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1279 = {{8'd0}, regs_1_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_700 = _T_698 - _GEN_1279; // @[Conwaylife.scala 29:42]
  wire  _T_701 = _T_700 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_702 = _T_700 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_703 = _T_700 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_705 = regs_1_15 + regs_1_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1280 = {{1'd0}, regs_1_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_706 = _T_705 + _GEN_1280; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1281 = {{2'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_707 = _T_706 + _GEN_1281; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1282 = {{3'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_708 = _T_707 + _GEN_1282; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1283 = {{4'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_709 = _T_708 + _GEN_1283; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1284 = {{5'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_710 = _T_709 + _GEN_1284; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1285 = {{6'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_711 = _T_710 + _GEN_1285; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1286 = {{7'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_712 = _T_711 + _GEN_1286; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1287 = {{8'd0}, regs_2_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_714 = _T_712 - _GEN_1287; // @[Conwaylife.scala 29:42]
  wire  _T_715 = _T_714 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_716 = _T_714 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_717 = _T_714 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_719 = regs_1_0 + regs_1_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1288 = {{1'd0}, regs_1_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_720 = _T_719 + _GEN_1288; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1289 = {{2'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_721 = _T_720 + _GEN_1289; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1290 = {{3'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_722 = _T_721 + _GEN_1290; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1291 = {{4'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_723 = _T_722 + _GEN_1291; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1292 = {{5'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_724 = _T_723 + _GEN_1292; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1293 = {{6'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_725 = _T_724 + _GEN_1293; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1294 = {{7'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_726 = _T_725 + _GEN_1294; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1295 = {{8'd0}, regs_2_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_728 = _T_726 - _GEN_1295; // @[Conwaylife.scala 29:42]
  wire  _T_729 = _T_728 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_730 = _T_728 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_731 = _T_728 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_733 = regs_1_1 + regs_1_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1296 = {{1'd0}, regs_1_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_734 = _T_733 + _GEN_1296; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1297 = {{2'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_735 = _T_734 + _GEN_1297; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1298 = {{3'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_736 = _T_735 + _GEN_1298; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1299 = {{4'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_737 = _T_736 + _GEN_1299; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1300 = {{5'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_738 = _T_737 + _GEN_1300; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1301 = {{6'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_739 = _T_738 + _GEN_1301; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1302 = {{7'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_740 = _T_739 + _GEN_1302; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1303 = {{8'd0}, regs_2_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_742 = _T_740 - _GEN_1303; // @[Conwaylife.scala 29:42]
  wire  _T_743 = _T_742 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_744 = _T_742 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_745 = _T_742 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_747 = regs_1_2 + regs_1_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1304 = {{1'd0}, regs_1_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_748 = _T_747 + _GEN_1304; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1305 = {{2'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_749 = _T_748 + _GEN_1305; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1306 = {{3'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_750 = _T_749 + _GEN_1306; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1307 = {{4'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_751 = _T_750 + _GEN_1307; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1308 = {{5'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_752 = _T_751 + _GEN_1308; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1309 = {{6'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_753 = _T_752 + _GEN_1309; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1310 = {{7'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_754 = _T_753 + _GEN_1310; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1311 = {{8'd0}, regs_2_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_756 = _T_754 - _GEN_1311; // @[Conwaylife.scala 29:42]
  wire  _T_757 = _T_756 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_758 = _T_756 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_759 = _T_756 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_761 = regs_1_3 + regs_1_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1312 = {{1'd0}, regs_1_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_762 = _T_761 + _GEN_1312; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1313 = {{2'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_763 = _T_762 + _GEN_1313; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1314 = {{3'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_764 = _T_763 + _GEN_1314; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1315 = {{4'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_765 = _T_764 + _GEN_1315; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1316 = {{5'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_766 = _T_765 + _GEN_1316; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1317 = {{6'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_767 = _T_766 + _GEN_1317; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1318 = {{7'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_768 = _T_767 + _GEN_1318; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1319 = {{8'd0}, regs_2_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_770 = _T_768 - _GEN_1319; // @[Conwaylife.scala 29:42]
  wire  _T_771 = _T_770 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_772 = _T_770 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_773 = _T_770 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_775 = regs_1_4 + regs_1_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1320 = {{1'd0}, regs_1_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_776 = _T_775 + _GEN_1320; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1321 = {{2'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_777 = _T_776 + _GEN_1321; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1322 = {{3'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_778 = _T_777 + _GEN_1322; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1323 = {{4'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_779 = _T_778 + _GEN_1323; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1324 = {{5'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_780 = _T_779 + _GEN_1324; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1325 = {{6'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_781 = _T_780 + _GEN_1325; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1326 = {{7'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_782 = _T_781 + _GEN_1326; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1327 = {{8'd0}, regs_2_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_784 = _T_782 - _GEN_1327; // @[Conwaylife.scala 29:42]
  wire  _T_785 = _T_784 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_786 = _T_784 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_787 = _T_784 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_789 = regs_1_5 + regs_1_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1328 = {{1'd0}, regs_1_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_790 = _T_789 + _GEN_1328; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1329 = {{2'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_791 = _T_790 + _GEN_1329; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1330 = {{3'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_792 = _T_791 + _GEN_1330; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1331 = {{4'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_793 = _T_792 + _GEN_1331; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1332 = {{5'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_794 = _T_793 + _GEN_1332; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1333 = {{6'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_795 = _T_794 + _GEN_1333; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1334 = {{7'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_796 = _T_795 + _GEN_1334; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1335 = {{8'd0}, regs_2_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_798 = _T_796 - _GEN_1335; // @[Conwaylife.scala 29:42]
  wire  _T_799 = _T_798 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_800 = _T_798 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_801 = _T_798 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_803 = regs_1_6 + regs_1_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1336 = {{1'd0}, regs_1_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_804 = _T_803 + _GEN_1336; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1337 = {{2'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_805 = _T_804 + _GEN_1337; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1338 = {{3'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_806 = _T_805 + _GEN_1338; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1339 = {{4'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_807 = _T_806 + _GEN_1339; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1340 = {{5'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_808 = _T_807 + _GEN_1340; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1341 = {{6'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_809 = _T_808 + _GEN_1341; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1342 = {{7'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_810 = _T_809 + _GEN_1342; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1343 = {{8'd0}, regs_2_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_812 = _T_810 - _GEN_1343; // @[Conwaylife.scala 29:42]
  wire  _T_813 = _T_812 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_814 = _T_812 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_815 = _T_812 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_817 = regs_1_7 + regs_1_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1344 = {{1'd0}, regs_1_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_818 = _T_817 + _GEN_1344; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1345 = {{2'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_819 = _T_818 + _GEN_1345; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1346 = {{3'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_820 = _T_819 + _GEN_1346; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1347 = {{4'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_821 = _T_820 + _GEN_1347; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1348 = {{5'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_822 = _T_821 + _GEN_1348; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1349 = {{6'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_823 = _T_822 + _GEN_1349; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1350 = {{7'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_824 = _T_823 + _GEN_1350; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1351 = {{8'd0}, regs_2_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_826 = _T_824 - _GEN_1351; // @[Conwaylife.scala 29:42]
  wire  _T_827 = _T_826 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_828 = _T_826 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_829 = _T_826 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_831 = regs_1_8 + regs_1_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1352 = {{1'd0}, regs_1_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_832 = _T_831 + _GEN_1352; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1353 = {{2'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_833 = _T_832 + _GEN_1353; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1354 = {{3'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_834 = _T_833 + _GEN_1354; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1355 = {{4'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_835 = _T_834 + _GEN_1355; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1356 = {{5'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_836 = _T_835 + _GEN_1356; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1357 = {{6'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_837 = _T_836 + _GEN_1357; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1358 = {{7'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_838 = _T_837 + _GEN_1358; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1359 = {{8'd0}, regs_2_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_840 = _T_838 - _GEN_1359; // @[Conwaylife.scala 29:42]
  wire  _T_841 = _T_840 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_842 = _T_840 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_843 = _T_840 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_845 = regs_1_9 + regs_1_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1360 = {{1'd0}, regs_1_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_846 = _T_845 + _GEN_1360; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1361 = {{2'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_847 = _T_846 + _GEN_1361; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1362 = {{3'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_848 = _T_847 + _GEN_1362; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1363 = {{4'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_849 = _T_848 + _GEN_1363; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1364 = {{5'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_850 = _T_849 + _GEN_1364; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1365 = {{6'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_851 = _T_850 + _GEN_1365; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1366 = {{7'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_852 = _T_851 + _GEN_1366; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1367 = {{8'd0}, regs_2_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_854 = _T_852 - _GEN_1367; // @[Conwaylife.scala 29:42]
  wire  _T_855 = _T_854 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_856 = _T_854 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_857 = _T_854 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_859 = regs_1_10 + regs_1_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1368 = {{1'd0}, regs_1_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_860 = _T_859 + _GEN_1368; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1369 = {{2'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_861 = _T_860 + _GEN_1369; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1370 = {{3'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_862 = _T_861 + _GEN_1370; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1371 = {{4'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_863 = _T_862 + _GEN_1371; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1372 = {{5'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_864 = _T_863 + _GEN_1372; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1373 = {{6'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_865 = _T_864 + _GEN_1373; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1374 = {{7'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_866 = _T_865 + _GEN_1374; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1375 = {{8'd0}, regs_2_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_868 = _T_866 - _GEN_1375; // @[Conwaylife.scala 29:42]
  wire  _T_869 = _T_868 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_870 = _T_868 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_871 = _T_868 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_873 = regs_1_11 + regs_1_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1376 = {{1'd0}, regs_1_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_874 = _T_873 + _GEN_1376; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1377 = {{2'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_875 = _T_874 + _GEN_1377; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1378 = {{3'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_876 = _T_875 + _GEN_1378; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1379 = {{4'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_877 = _T_876 + _GEN_1379; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1380 = {{5'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_878 = _T_877 + _GEN_1380; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1381 = {{6'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_879 = _T_878 + _GEN_1381; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1382 = {{7'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_880 = _T_879 + _GEN_1382; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1383 = {{8'd0}, regs_2_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_882 = _T_880 - _GEN_1383; // @[Conwaylife.scala 29:42]
  wire  _T_883 = _T_882 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_884 = _T_882 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_885 = _T_882 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_887 = regs_1_12 + regs_1_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1384 = {{1'd0}, regs_1_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_888 = _T_887 + _GEN_1384; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1385 = {{2'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_889 = _T_888 + _GEN_1385; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1386 = {{3'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_890 = _T_889 + _GEN_1386; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1387 = {{4'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_891 = _T_890 + _GEN_1387; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1388 = {{5'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_892 = _T_891 + _GEN_1388; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1389 = {{6'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_893 = _T_892 + _GEN_1389; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1390 = {{7'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_894 = _T_893 + _GEN_1390; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1391 = {{8'd0}, regs_2_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_896 = _T_894 - _GEN_1391; // @[Conwaylife.scala 29:42]
  wire  _T_897 = _T_896 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_898 = _T_896 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_899 = _T_896 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_901 = regs_1_13 + regs_1_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1392 = {{1'd0}, regs_1_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_902 = _T_901 + _GEN_1392; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1393 = {{2'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_903 = _T_902 + _GEN_1393; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1394 = {{3'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_904 = _T_903 + _GEN_1394; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1395 = {{4'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_905 = _T_904 + _GEN_1395; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1396 = {{5'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_906 = _T_905 + _GEN_1396; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1397 = {{6'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_907 = _T_906 + _GEN_1397; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1398 = {{7'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_908 = _T_907 + _GEN_1398; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1399 = {{8'd0}, regs_2_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_910 = _T_908 - _GEN_1399; // @[Conwaylife.scala 29:42]
  wire  _T_911 = _T_910 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_912 = _T_910 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_913 = _T_910 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_915 = regs_1_14 + regs_1_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1400 = {{1'd0}, regs_1_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_916 = _T_915 + _GEN_1400; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1401 = {{2'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_917 = _T_916 + _GEN_1401; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1402 = {{3'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_918 = _T_917 + _GEN_1402; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1403 = {{4'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_919 = _T_918 + _GEN_1403; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1404 = {{5'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_920 = _T_919 + _GEN_1404; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1405 = {{6'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_921 = _T_920 + _GEN_1405; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1406 = {{7'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_922 = _T_921 + _GEN_1406; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1407 = {{8'd0}, regs_2_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_924 = _T_922 - _GEN_1407; // @[Conwaylife.scala 29:42]
  wire  _T_925 = _T_924 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_926 = _T_924 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_927 = _T_924 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_929 = regs_2_15 + regs_2_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1408 = {{1'd0}, regs_2_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_930 = _T_929 + _GEN_1408; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1409 = {{2'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_931 = _T_930 + _GEN_1409; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1410 = {{3'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_932 = _T_931 + _GEN_1410; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1411 = {{4'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_933 = _T_932 + _GEN_1411; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1412 = {{5'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_934 = _T_933 + _GEN_1412; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1413 = {{6'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_935 = _T_934 + _GEN_1413; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1414 = {{7'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_936 = _T_935 + _GEN_1414; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1415 = {{8'd0}, regs_3_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_938 = _T_936 - _GEN_1415; // @[Conwaylife.scala 29:42]
  wire  _T_939 = _T_938 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_940 = _T_938 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_941 = _T_938 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_943 = regs_2_0 + regs_2_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1416 = {{1'd0}, regs_2_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_944 = _T_943 + _GEN_1416; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1417 = {{2'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_945 = _T_944 + _GEN_1417; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1418 = {{3'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_946 = _T_945 + _GEN_1418; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1419 = {{4'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_947 = _T_946 + _GEN_1419; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1420 = {{5'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_948 = _T_947 + _GEN_1420; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1421 = {{6'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_949 = _T_948 + _GEN_1421; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1422 = {{7'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_950 = _T_949 + _GEN_1422; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1423 = {{8'd0}, regs_3_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_952 = _T_950 - _GEN_1423; // @[Conwaylife.scala 29:42]
  wire  _T_953 = _T_952 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_954 = _T_952 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_955 = _T_952 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_957 = regs_2_1 + regs_2_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1424 = {{1'd0}, regs_2_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_958 = _T_957 + _GEN_1424; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1425 = {{2'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_959 = _T_958 + _GEN_1425; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1426 = {{3'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_960 = _T_959 + _GEN_1426; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1427 = {{4'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_961 = _T_960 + _GEN_1427; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1428 = {{5'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_962 = _T_961 + _GEN_1428; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1429 = {{6'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_963 = _T_962 + _GEN_1429; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1430 = {{7'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_964 = _T_963 + _GEN_1430; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1431 = {{8'd0}, regs_3_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_966 = _T_964 - _GEN_1431; // @[Conwaylife.scala 29:42]
  wire  _T_967 = _T_966 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_968 = _T_966 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_969 = _T_966 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_971 = regs_2_2 + regs_2_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1432 = {{1'd0}, regs_2_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_972 = _T_971 + _GEN_1432; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1433 = {{2'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_973 = _T_972 + _GEN_1433; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1434 = {{3'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_974 = _T_973 + _GEN_1434; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1435 = {{4'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_975 = _T_974 + _GEN_1435; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1436 = {{5'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_976 = _T_975 + _GEN_1436; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1437 = {{6'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_977 = _T_976 + _GEN_1437; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1438 = {{7'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_978 = _T_977 + _GEN_1438; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1439 = {{8'd0}, regs_3_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_980 = _T_978 - _GEN_1439; // @[Conwaylife.scala 29:42]
  wire  _T_981 = _T_980 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_982 = _T_980 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_983 = _T_980 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_985 = regs_2_3 + regs_2_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1440 = {{1'd0}, regs_2_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_986 = _T_985 + _GEN_1440; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1441 = {{2'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_987 = _T_986 + _GEN_1441; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1442 = {{3'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_988 = _T_987 + _GEN_1442; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1443 = {{4'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_989 = _T_988 + _GEN_1443; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1444 = {{5'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_990 = _T_989 + _GEN_1444; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1445 = {{6'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_991 = _T_990 + _GEN_1445; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1446 = {{7'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_992 = _T_991 + _GEN_1446; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1447 = {{8'd0}, regs_3_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_994 = _T_992 - _GEN_1447; // @[Conwaylife.scala 29:42]
  wire  _T_995 = _T_994 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_996 = _T_994 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_997 = _T_994 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_999 = regs_2_4 + regs_2_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1448 = {{1'd0}, regs_2_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1000 = _T_999 + _GEN_1448; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1449 = {{2'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1001 = _T_1000 + _GEN_1449; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1450 = {{3'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1002 = _T_1001 + _GEN_1450; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1451 = {{4'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1003 = _T_1002 + _GEN_1451; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1452 = {{5'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1004 = _T_1003 + _GEN_1452; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1453 = {{6'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1005 = _T_1004 + _GEN_1453; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1454 = {{7'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1006 = _T_1005 + _GEN_1454; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1455 = {{8'd0}, regs_3_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1008 = _T_1006 - _GEN_1455; // @[Conwaylife.scala 29:42]
  wire  _T_1009 = _T_1008 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1010 = _T_1008 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1011 = _T_1008 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1013 = regs_2_5 + regs_2_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1456 = {{1'd0}, regs_2_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1014 = _T_1013 + _GEN_1456; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1457 = {{2'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1015 = _T_1014 + _GEN_1457; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1458 = {{3'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1016 = _T_1015 + _GEN_1458; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1459 = {{4'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1017 = _T_1016 + _GEN_1459; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1460 = {{5'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1018 = _T_1017 + _GEN_1460; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1461 = {{6'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1019 = _T_1018 + _GEN_1461; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1462 = {{7'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1020 = _T_1019 + _GEN_1462; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1463 = {{8'd0}, regs_3_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1022 = _T_1020 - _GEN_1463; // @[Conwaylife.scala 29:42]
  wire  _T_1023 = _T_1022 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1024 = _T_1022 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1025 = _T_1022 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1027 = regs_2_6 + regs_2_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1464 = {{1'd0}, regs_2_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1028 = _T_1027 + _GEN_1464; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1465 = {{2'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1029 = _T_1028 + _GEN_1465; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1466 = {{3'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1030 = _T_1029 + _GEN_1466; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1467 = {{4'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1031 = _T_1030 + _GEN_1467; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1468 = {{5'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1032 = _T_1031 + _GEN_1468; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1469 = {{6'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1033 = _T_1032 + _GEN_1469; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1470 = {{7'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1034 = _T_1033 + _GEN_1470; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1471 = {{8'd0}, regs_3_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1036 = _T_1034 - _GEN_1471; // @[Conwaylife.scala 29:42]
  wire  _T_1037 = _T_1036 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1038 = _T_1036 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1039 = _T_1036 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1041 = regs_2_7 + regs_2_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1472 = {{1'd0}, regs_2_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1042 = _T_1041 + _GEN_1472; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1473 = {{2'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1043 = _T_1042 + _GEN_1473; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1474 = {{3'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1044 = _T_1043 + _GEN_1474; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1475 = {{4'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1045 = _T_1044 + _GEN_1475; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1476 = {{5'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1046 = _T_1045 + _GEN_1476; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1477 = {{6'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1047 = _T_1046 + _GEN_1477; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1478 = {{7'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1048 = _T_1047 + _GEN_1478; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1479 = {{8'd0}, regs_3_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1050 = _T_1048 - _GEN_1479; // @[Conwaylife.scala 29:42]
  wire  _T_1051 = _T_1050 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1052 = _T_1050 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1053 = _T_1050 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1055 = regs_2_8 + regs_2_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1480 = {{1'd0}, regs_2_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1056 = _T_1055 + _GEN_1480; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1481 = {{2'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1057 = _T_1056 + _GEN_1481; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1482 = {{3'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1058 = _T_1057 + _GEN_1482; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1483 = {{4'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1059 = _T_1058 + _GEN_1483; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1484 = {{5'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1060 = _T_1059 + _GEN_1484; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1485 = {{6'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1061 = _T_1060 + _GEN_1485; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1486 = {{7'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1062 = _T_1061 + _GEN_1486; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1487 = {{8'd0}, regs_3_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1064 = _T_1062 - _GEN_1487; // @[Conwaylife.scala 29:42]
  wire  _T_1065 = _T_1064 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1066 = _T_1064 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1067 = _T_1064 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1069 = regs_2_9 + regs_2_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1488 = {{1'd0}, regs_2_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1070 = _T_1069 + _GEN_1488; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1489 = {{2'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1071 = _T_1070 + _GEN_1489; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1490 = {{3'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1072 = _T_1071 + _GEN_1490; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1491 = {{4'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1073 = _T_1072 + _GEN_1491; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1492 = {{5'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1074 = _T_1073 + _GEN_1492; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1493 = {{6'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1075 = _T_1074 + _GEN_1493; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1494 = {{7'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1076 = _T_1075 + _GEN_1494; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1495 = {{8'd0}, regs_3_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1078 = _T_1076 - _GEN_1495; // @[Conwaylife.scala 29:42]
  wire  _T_1079 = _T_1078 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1080 = _T_1078 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1081 = _T_1078 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1083 = regs_2_10 + regs_2_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1496 = {{1'd0}, regs_2_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1084 = _T_1083 + _GEN_1496; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1497 = {{2'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1085 = _T_1084 + _GEN_1497; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1498 = {{3'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1086 = _T_1085 + _GEN_1498; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1499 = {{4'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1087 = _T_1086 + _GEN_1499; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1500 = {{5'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1088 = _T_1087 + _GEN_1500; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1501 = {{6'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1089 = _T_1088 + _GEN_1501; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1502 = {{7'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1090 = _T_1089 + _GEN_1502; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1503 = {{8'd0}, regs_3_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1092 = _T_1090 - _GEN_1503; // @[Conwaylife.scala 29:42]
  wire  _T_1093 = _T_1092 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1094 = _T_1092 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1095 = _T_1092 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1097 = regs_2_11 + regs_2_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1504 = {{1'd0}, regs_2_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1098 = _T_1097 + _GEN_1504; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1505 = {{2'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1099 = _T_1098 + _GEN_1505; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1506 = {{3'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1100 = _T_1099 + _GEN_1506; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1507 = {{4'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1101 = _T_1100 + _GEN_1507; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1508 = {{5'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1102 = _T_1101 + _GEN_1508; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1509 = {{6'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1103 = _T_1102 + _GEN_1509; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1510 = {{7'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1104 = _T_1103 + _GEN_1510; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1511 = {{8'd0}, regs_3_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1106 = _T_1104 - _GEN_1511; // @[Conwaylife.scala 29:42]
  wire  _T_1107 = _T_1106 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1108 = _T_1106 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1109 = _T_1106 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1111 = regs_2_12 + regs_2_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1512 = {{1'd0}, regs_2_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1112 = _T_1111 + _GEN_1512; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1513 = {{2'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1113 = _T_1112 + _GEN_1513; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1514 = {{3'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1114 = _T_1113 + _GEN_1514; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1515 = {{4'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1115 = _T_1114 + _GEN_1515; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1516 = {{5'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1116 = _T_1115 + _GEN_1516; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1517 = {{6'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1117 = _T_1116 + _GEN_1517; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1518 = {{7'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1118 = _T_1117 + _GEN_1518; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1519 = {{8'd0}, regs_3_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1120 = _T_1118 - _GEN_1519; // @[Conwaylife.scala 29:42]
  wire  _T_1121 = _T_1120 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1122 = _T_1120 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1123 = _T_1120 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1125 = regs_2_13 + regs_2_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1520 = {{1'd0}, regs_2_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1126 = _T_1125 + _GEN_1520; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1521 = {{2'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1127 = _T_1126 + _GEN_1521; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1522 = {{3'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1128 = _T_1127 + _GEN_1522; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1523 = {{4'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1129 = _T_1128 + _GEN_1523; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1524 = {{5'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1130 = _T_1129 + _GEN_1524; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1525 = {{6'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1131 = _T_1130 + _GEN_1525; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1526 = {{7'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1132 = _T_1131 + _GEN_1526; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1527 = {{8'd0}, regs_3_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1134 = _T_1132 - _GEN_1527; // @[Conwaylife.scala 29:42]
  wire  _T_1135 = _T_1134 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1136 = _T_1134 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1137 = _T_1134 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1139 = regs_2_14 + regs_2_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1528 = {{1'd0}, regs_2_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1140 = _T_1139 + _GEN_1528; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1529 = {{2'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1141 = _T_1140 + _GEN_1529; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1530 = {{3'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1142 = _T_1141 + _GEN_1530; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1531 = {{4'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1143 = _T_1142 + _GEN_1531; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1532 = {{5'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1144 = _T_1143 + _GEN_1532; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1533 = {{6'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1145 = _T_1144 + _GEN_1533; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1534 = {{7'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1146 = _T_1145 + _GEN_1534; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1535 = {{8'd0}, regs_3_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1148 = _T_1146 - _GEN_1535; // @[Conwaylife.scala 29:42]
  wire  _T_1149 = _T_1148 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1150 = _T_1148 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1151 = _T_1148 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1153 = regs_3_15 + regs_3_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1536 = {{1'd0}, regs_3_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1154 = _T_1153 + _GEN_1536; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1537 = {{2'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1155 = _T_1154 + _GEN_1537; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1538 = {{3'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1156 = _T_1155 + _GEN_1538; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1539 = {{4'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1157 = _T_1156 + _GEN_1539; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1540 = {{5'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1158 = _T_1157 + _GEN_1540; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1541 = {{6'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1159 = _T_1158 + _GEN_1541; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1542 = {{7'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1160 = _T_1159 + _GEN_1542; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1543 = {{8'd0}, regs_4_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1162 = _T_1160 - _GEN_1543; // @[Conwaylife.scala 29:42]
  wire  _T_1163 = _T_1162 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1164 = _T_1162 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1165 = _T_1162 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1167 = regs_3_0 + regs_3_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1544 = {{1'd0}, regs_3_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1168 = _T_1167 + _GEN_1544; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1545 = {{2'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1169 = _T_1168 + _GEN_1545; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1546 = {{3'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1170 = _T_1169 + _GEN_1546; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1547 = {{4'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1171 = _T_1170 + _GEN_1547; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1548 = {{5'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1172 = _T_1171 + _GEN_1548; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1549 = {{6'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1173 = _T_1172 + _GEN_1549; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1550 = {{7'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1174 = _T_1173 + _GEN_1550; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1551 = {{8'd0}, regs_4_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1176 = _T_1174 - _GEN_1551; // @[Conwaylife.scala 29:42]
  wire  _T_1177 = _T_1176 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1178 = _T_1176 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1179 = _T_1176 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1181 = regs_3_1 + regs_3_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1552 = {{1'd0}, regs_3_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1182 = _T_1181 + _GEN_1552; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1553 = {{2'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1183 = _T_1182 + _GEN_1553; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1554 = {{3'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1184 = _T_1183 + _GEN_1554; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1555 = {{4'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1185 = _T_1184 + _GEN_1555; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1556 = {{5'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1186 = _T_1185 + _GEN_1556; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1557 = {{6'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1187 = _T_1186 + _GEN_1557; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1558 = {{7'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1188 = _T_1187 + _GEN_1558; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1559 = {{8'd0}, regs_4_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1190 = _T_1188 - _GEN_1559; // @[Conwaylife.scala 29:42]
  wire  _T_1191 = _T_1190 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1192 = _T_1190 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1193 = _T_1190 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1195 = regs_3_2 + regs_3_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1560 = {{1'd0}, regs_3_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1196 = _T_1195 + _GEN_1560; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1561 = {{2'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1197 = _T_1196 + _GEN_1561; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1562 = {{3'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1198 = _T_1197 + _GEN_1562; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1563 = {{4'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1199 = _T_1198 + _GEN_1563; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1564 = {{5'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1200 = _T_1199 + _GEN_1564; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1565 = {{6'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1201 = _T_1200 + _GEN_1565; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1566 = {{7'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1202 = _T_1201 + _GEN_1566; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1567 = {{8'd0}, regs_4_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1204 = _T_1202 - _GEN_1567; // @[Conwaylife.scala 29:42]
  wire  _T_1205 = _T_1204 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1206 = _T_1204 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1207 = _T_1204 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1209 = regs_3_3 + regs_3_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1568 = {{1'd0}, regs_3_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1210 = _T_1209 + _GEN_1568; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1569 = {{2'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1211 = _T_1210 + _GEN_1569; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1570 = {{3'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1212 = _T_1211 + _GEN_1570; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1571 = {{4'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1213 = _T_1212 + _GEN_1571; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1572 = {{5'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1214 = _T_1213 + _GEN_1572; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1573 = {{6'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1215 = _T_1214 + _GEN_1573; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1574 = {{7'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1216 = _T_1215 + _GEN_1574; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1575 = {{8'd0}, regs_4_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1218 = _T_1216 - _GEN_1575; // @[Conwaylife.scala 29:42]
  wire  _T_1219 = _T_1218 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1220 = _T_1218 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1221 = _T_1218 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1223 = regs_3_4 + regs_3_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1576 = {{1'd0}, regs_3_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1224 = _T_1223 + _GEN_1576; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1577 = {{2'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1225 = _T_1224 + _GEN_1577; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1578 = {{3'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1226 = _T_1225 + _GEN_1578; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1579 = {{4'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1227 = _T_1226 + _GEN_1579; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1580 = {{5'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1228 = _T_1227 + _GEN_1580; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1581 = {{6'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1229 = _T_1228 + _GEN_1581; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1582 = {{7'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1230 = _T_1229 + _GEN_1582; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1583 = {{8'd0}, regs_4_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1232 = _T_1230 - _GEN_1583; // @[Conwaylife.scala 29:42]
  wire  _T_1233 = _T_1232 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1234 = _T_1232 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1235 = _T_1232 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1237 = regs_3_5 + regs_3_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1584 = {{1'd0}, regs_3_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1238 = _T_1237 + _GEN_1584; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1585 = {{2'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1239 = _T_1238 + _GEN_1585; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1586 = {{3'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1240 = _T_1239 + _GEN_1586; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1587 = {{4'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1241 = _T_1240 + _GEN_1587; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1588 = {{5'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1242 = _T_1241 + _GEN_1588; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1589 = {{6'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1243 = _T_1242 + _GEN_1589; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1590 = {{7'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1244 = _T_1243 + _GEN_1590; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1591 = {{8'd0}, regs_4_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1246 = _T_1244 - _GEN_1591; // @[Conwaylife.scala 29:42]
  wire  _T_1247 = _T_1246 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1248 = _T_1246 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1249 = _T_1246 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1251 = regs_3_6 + regs_3_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1592 = {{1'd0}, regs_3_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1252 = _T_1251 + _GEN_1592; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1593 = {{2'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1253 = _T_1252 + _GEN_1593; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1594 = {{3'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1254 = _T_1253 + _GEN_1594; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1595 = {{4'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1255 = _T_1254 + _GEN_1595; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1596 = {{5'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1256 = _T_1255 + _GEN_1596; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1597 = {{6'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1257 = _T_1256 + _GEN_1597; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1598 = {{7'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1258 = _T_1257 + _GEN_1598; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1599 = {{8'd0}, regs_4_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1260 = _T_1258 - _GEN_1599; // @[Conwaylife.scala 29:42]
  wire  _T_1261 = _T_1260 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1262 = _T_1260 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1263 = _T_1260 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1265 = regs_3_7 + regs_3_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1600 = {{1'd0}, regs_3_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1266 = _T_1265 + _GEN_1600; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1601 = {{2'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1267 = _T_1266 + _GEN_1601; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1602 = {{3'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1268 = _T_1267 + _GEN_1602; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1603 = {{4'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1269 = _T_1268 + _GEN_1603; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1604 = {{5'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1270 = _T_1269 + _GEN_1604; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1605 = {{6'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1271 = _T_1270 + _GEN_1605; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1606 = {{7'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1272 = _T_1271 + _GEN_1606; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1607 = {{8'd0}, regs_4_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1274 = _T_1272 - _GEN_1607; // @[Conwaylife.scala 29:42]
  wire  _T_1275 = _T_1274 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1276 = _T_1274 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1277 = _T_1274 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1279 = regs_3_8 + regs_3_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1608 = {{1'd0}, regs_3_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1280 = _T_1279 + _GEN_1608; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1609 = {{2'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1281 = _T_1280 + _GEN_1609; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1610 = {{3'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1282 = _T_1281 + _GEN_1610; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1611 = {{4'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1283 = _T_1282 + _GEN_1611; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1612 = {{5'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1284 = _T_1283 + _GEN_1612; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1613 = {{6'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1285 = _T_1284 + _GEN_1613; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1614 = {{7'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1286 = _T_1285 + _GEN_1614; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1615 = {{8'd0}, regs_4_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1288 = _T_1286 - _GEN_1615; // @[Conwaylife.scala 29:42]
  wire  _T_1289 = _T_1288 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1290 = _T_1288 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1291 = _T_1288 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1293 = regs_3_9 + regs_3_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1616 = {{1'd0}, regs_3_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1294 = _T_1293 + _GEN_1616; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1617 = {{2'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1295 = _T_1294 + _GEN_1617; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1618 = {{3'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1296 = _T_1295 + _GEN_1618; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1619 = {{4'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1297 = _T_1296 + _GEN_1619; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1620 = {{5'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1298 = _T_1297 + _GEN_1620; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1621 = {{6'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1299 = _T_1298 + _GEN_1621; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1622 = {{7'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1300 = _T_1299 + _GEN_1622; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1623 = {{8'd0}, regs_4_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1302 = _T_1300 - _GEN_1623; // @[Conwaylife.scala 29:42]
  wire  _T_1303 = _T_1302 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1304 = _T_1302 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1305 = _T_1302 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1307 = regs_3_10 + regs_3_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1624 = {{1'd0}, regs_3_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1308 = _T_1307 + _GEN_1624; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1625 = {{2'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1309 = _T_1308 + _GEN_1625; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1626 = {{3'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1310 = _T_1309 + _GEN_1626; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1627 = {{4'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1311 = _T_1310 + _GEN_1627; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1628 = {{5'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1312 = _T_1311 + _GEN_1628; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1629 = {{6'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1313 = _T_1312 + _GEN_1629; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1630 = {{7'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1314 = _T_1313 + _GEN_1630; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1631 = {{8'd0}, regs_4_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1316 = _T_1314 - _GEN_1631; // @[Conwaylife.scala 29:42]
  wire  _T_1317 = _T_1316 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1318 = _T_1316 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1319 = _T_1316 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1321 = regs_3_11 + regs_3_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1632 = {{1'd0}, regs_3_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1322 = _T_1321 + _GEN_1632; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1633 = {{2'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1323 = _T_1322 + _GEN_1633; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1634 = {{3'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1324 = _T_1323 + _GEN_1634; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1635 = {{4'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1325 = _T_1324 + _GEN_1635; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1636 = {{5'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1326 = _T_1325 + _GEN_1636; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1637 = {{6'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1327 = _T_1326 + _GEN_1637; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1638 = {{7'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1328 = _T_1327 + _GEN_1638; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1639 = {{8'd0}, regs_4_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1330 = _T_1328 - _GEN_1639; // @[Conwaylife.scala 29:42]
  wire  _T_1331 = _T_1330 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1332 = _T_1330 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1333 = _T_1330 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1335 = regs_3_12 + regs_3_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1640 = {{1'd0}, regs_3_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1336 = _T_1335 + _GEN_1640; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1641 = {{2'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1337 = _T_1336 + _GEN_1641; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1642 = {{3'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1338 = _T_1337 + _GEN_1642; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1643 = {{4'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1339 = _T_1338 + _GEN_1643; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1644 = {{5'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1340 = _T_1339 + _GEN_1644; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1645 = {{6'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1341 = _T_1340 + _GEN_1645; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1646 = {{7'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1342 = _T_1341 + _GEN_1646; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1647 = {{8'd0}, regs_4_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1344 = _T_1342 - _GEN_1647; // @[Conwaylife.scala 29:42]
  wire  _T_1345 = _T_1344 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1346 = _T_1344 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1347 = _T_1344 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1349 = regs_3_13 + regs_3_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1648 = {{1'd0}, regs_3_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1350 = _T_1349 + _GEN_1648; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1649 = {{2'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1351 = _T_1350 + _GEN_1649; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1650 = {{3'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1352 = _T_1351 + _GEN_1650; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1651 = {{4'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1353 = _T_1352 + _GEN_1651; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1652 = {{5'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1354 = _T_1353 + _GEN_1652; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1653 = {{6'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1355 = _T_1354 + _GEN_1653; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1654 = {{7'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1356 = _T_1355 + _GEN_1654; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1655 = {{8'd0}, regs_4_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1358 = _T_1356 - _GEN_1655; // @[Conwaylife.scala 29:42]
  wire  _T_1359 = _T_1358 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1360 = _T_1358 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1361 = _T_1358 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1363 = regs_3_14 + regs_3_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1656 = {{1'd0}, regs_3_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1364 = _T_1363 + _GEN_1656; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1657 = {{2'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1365 = _T_1364 + _GEN_1657; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1658 = {{3'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1366 = _T_1365 + _GEN_1658; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1659 = {{4'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1367 = _T_1366 + _GEN_1659; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1660 = {{5'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1368 = _T_1367 + _GEN_1660; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1661 = {{6'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1369 = _T_1368 + _GEN_1661; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1662 = {{7'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1370 = _T_1369 + _GEN_1662; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1663 = {{8'd0}, regs_4_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1372 = _T_1370 - _GEN_1663; // @[Conwaylife.scala 29:42]
  wire  _T_1373 = _T_1372 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1374 = _T_1372 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1375 = _T_1372 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1377 = regs_4_15 + regs_4_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1664 = {{1'd0}, regs_4_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1378 = _T_1377 + _GEN_1664; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1665 = {{2'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1379 = _T_1378 + _GEN_1665; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1666 = {{3'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1380 = _T_1379 + _GEN_1666; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1667 = {{4'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1381 = _T_1380 + _GEN_1667; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1668 = {{5'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1382 = _T_1381 + _GEN_1668; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1669 = {{6'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1383 = _T_1382 + _GEN_1669; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1670 = {{7'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1384 = _T_1383 + _GEN_1670; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1671 = {{8'd0}, regs_5_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1386 = _T_1384 - _GEN_1671; // @[Conwaylife.scala 29:42]
  wire  _T_1387 = _T_1386 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1388 = _T_1386 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1389 = _T_1386 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1391 = regs_4_0 + regs_4_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1672 = {{1'd0}, regs_4_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1392 = _T_1391 + _GEN_1672; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1673 = {{2'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1393 = _T_1392 + _GEN_1673; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1674 = {{3'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1394 = _T_1393 + _GEN_1674; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1675 = {{4'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1395 = _T_1394 + _GEN_1675; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1676 = {{5'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1396 = _T_1395 + _GEN_1676; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1677 = {{6'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1397 = _T_1396 + _GEN_1677; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1678 = {{7'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1398 = _T_1397 + _GEN_1678; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1679 = {{8'd0}, regs_5_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1400 = _T_1398 - _GEN_1679; // @[Conwaylife.scala 29:42]
  wire  _T_1401 = _T_1400 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1402 = _T_1400 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1403 = _T_1400 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1405 = regs_4_1 + regs_4_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1680 = {{1'd0}, regs_4_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1406 = _T_1405 + _GEN_1680; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1681 = {{2'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1407 = _T_1406 + _GEN_1681; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1682 = {{3'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1408 = _T_1407 + _GEN_1682; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1683 = {{4'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1409 = _T_1408 + _GEN_1683; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1684 = {{5'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1410 = _T_1409 + _GEN_1684; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1685 = {{6'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1411 = _T_1410 + _GEN_1685; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1686 = {{7'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1412 = _T_1411 + _GEN_1686; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1687 = {{8'd0}, regs_5_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1414 = _T_1412 - _GEN_1687; // @[Conwaylife.scala 29:42]
  wire  _T_1415 = _T_1414 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1416 = _T_1414 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1417 = _T_1414 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1419 = regs_4_2 + regs_4_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1688 = {{1'd0}, regs_4_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1420 = _T_1419 + _GEN_1688; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1689 = {{2'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1421 = _T_1420 + _GEN_1689; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1690 = {{3'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1422 = _T_1421 + _GEN_1690; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1691 = {{4'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1423 = _T_1422 + _GEN_1691; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1692 = {{5'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1424 = _T_1423 + _GEN_1692; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1693 = {{6'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1425 = _T_1424 + _GEN_1693; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1694 = {{7'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1426 = _T_1425 + _GEN_1694; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1695 = {{8'd0}, regs_5_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1428 = _T_1426 - _GEN_1695; // @[Conwaylife.scala 29:42]
  wire  _T_1429 = _T_1428 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1430 = _T_1428 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1431 = _T_1428 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1433 = regs_4_3 + regs_4_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1696 = {{1'd0}, regs_4_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1434 = _T_1433 + _GEN_1696; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1697 = {{2'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1435 = _T_1434 + _GEN_1697; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1698 = {{3'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1436 = _T_1435 + _GEN_1698; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1699 = {{4'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1437 = _T_1436 + _GEN_1699; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1700 = {{5'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1438 = _T_1437 + _GEN_1700; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1701 = {{6'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1439 = _T_1438 + _GEN_1701; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1702 = {{7'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1440 = _T_1439 + _GEN_1702; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1703 = {{8'd0}, regs_5_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1442 = _T_1440 - _GEN_1703; // @[Conwaylife.scala 29:42]
  wire  _T_1443 = _T_1442 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1444 = _T_1442 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1445 = _T_1442 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1447 = regs_4_4 + regs_4_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1704 = {{1'd0}, regs_4_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1448 = _T_1447 + _GEN_1704; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1705 = {{2'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1449 = _T_1448 + _GEN_1705; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1706 = {{3'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1450 = _T_1449 + _GEN_1706; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1707 = {{4'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1451 = _T_1450 + _GEN_1707; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1708 = {{5'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1452 = _T_1451 + _GEN_1708; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1709 = {{6'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1453 = _T_1452 + _GEN_1709; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1710 = {{7'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1454 = _T_1453 + _GEN_1710; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1711 = {{8'd0}, regs_5_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1456 = _T_1454 - _GEN_1711; // @[Conwaylife.scala 29:42]
  wire  _T_1457 = _T_1456 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1458 = _T_1456 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1459 = _T_1456 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1461 = regs_4_5 + regs_4_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1712 = {{1'd0}, regs_4_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1462 = _T_1461 + _GEN_1712; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1713 = {{2'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1463 = _T_1462 + _GEN_1713; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1714 = {{3'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1464 = _T_1463 + _GEN_1714; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1715 = {{4'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1465 = _T_1464 + _GEN_1715; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1716 = {{5'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1466 = _T_1465 + _GEN_1716; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1717 = {{6'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1467 = _T_1466 + _GEN_1717; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1718 = {{7'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1468 = _T_1467 + _GEN_1718; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1719 = {{8'd0}, regs_5_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1470 = _T_1468 - _GEN_1719; // @[Conwaylife.scala 29:42]
  wire  _T_1471 = _T_1470 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1472 = _T_1470 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1473 = _T_1470 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1475 = regs_4_6 + regs_4_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1720 = {{1'd0}, regs_4_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1476 = _T_1475 + _GEN_1720; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1721 = {{2'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1477 = _T_1476 + _GEN_1721; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1722 = {{3'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1478 = _T_1477 + _GEN_1722; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1723 = {{4'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1479 = _T_1478 + _GEN_1723; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1724 = {{5'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1480 = _T_1479 + _GEN_1724; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1725 = {{6'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1481 = _T_1480 + _GEN_1725; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1726 = {{7'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1482 = _T_1481 + _GEN_1726; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1727 = {{8'd0}, regs_5_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1484 = _T_1482 - _GEN_1727; // @[Conwaylife.scala 29:42]
  wire  _T_1485 = _T_1484 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1486 = _T_1484 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1487 = _T_1484 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1489 = regs_4_7 + regs_4_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1728 = {{1'd0}, regs_4_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1490 = _T_1489 + _GEN_1728; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1729 = {{2'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1491 = _T_1490 + _GEN_1729; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1730 = {{3'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1492 = _T_1491 + _GEN_1730; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1731 = {{4'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1493 = _T_1492 + _GEN_1731; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1732 = {{5'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1494 = _T_1493 + _GEN_1732; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1733 = {{6'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1495 = _T_1494 + _GEN_1733; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1734 = {{7'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1496 = _T_1495 + _GEN_1734; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1735 = {{8'd0}, regs_5_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1498 = _T_1496 - _GEN_1735; // @[Conwaylife.scala 29:42]
  wire  _T_1499 = _T_1498 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1500 = _T_1498 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1501 = _T_1498 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1503 = regs_4_8 + regs_4_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1736 = {{1'd0}, regs_4_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1504 = _T_1503 + _GEN_1736; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1737 = {{2'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1505 = _T_1504 + _GEN_1737; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1738 = {{3'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1506 = _T_1505 + _GEN_1738; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1739 = {{4'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1507 = _T_1506 + _GEN_1739; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1740 = {{5'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1508 = _T_1507 + _GEN_1740; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1741 = {{6'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1509 = _T_1508 + _GEN_1741; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1742 = {{7'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1510 = _T_1509 + _GEN_1742; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1743 = {{8'd0}, regs_5_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1512 = _T_1510 - _GEN_1743; // @[Conwaylife.scala 29:42]
  wire  _T_1513 = _T_1512 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1514 = _T_1512 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1515 = _T_1512 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1517 = regs_4_9 + regs_4_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1744 = {{1'd0}, regs_4_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1518 = _T_1517 + _GEN_1744; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1745 = {{2'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1519 = _T_1518 + _GEN_1745; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1746 = {{3'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1520 = _T_1519 + _GEN_1746; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1747 = {{4'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1521 = _T_1520 + _GEN_1747; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1748 = {{5'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1522 = _T_1521 + _GEN_1748; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1749 = {{6'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1523 = _T_1522 + _GEN_1749; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1750 = {{7'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1524 = _T_1523 + _GEN_1750; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1751 = {{8'd0}, regs_5_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1526 = _T_1524 - _GEN_1751; // @[Conwaylife.scala 29:42]
  wire  _T_1527 = _T_1526 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1528 = _T_1526 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1529 = _T_1526 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1531 = regs_4_10 + regs_4_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1752 = {{1'd0}, regs_4_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1532 = _T_1531 + _GEN_1752; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1753 = {{2'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1533 = _T_1532 + _GEN_1753; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1754 = {{3'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1534 = _T_1533 + _GEN_1754; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1755 = {{4'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1535 = _T_1534 + _GEN_1755; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1756 = {{5'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1536 = _T_1535 + _GEN_1756; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1757 = {{6'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1537 = _T_1536 + _GEN_1757; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1758 = {{7'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1538 = _T_1537 + _GEN_1758; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1759 = {{8'd0}, regs_5_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1540 = _T_1538 - _GEN_1759; // @[Conwaylife.scala 29:42]
  wire  _T_1541 = _T_1540 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1542 = _T_1540 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1543 = _T_1540 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1545 = regs_4_11 + regs_4_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1760 = {{1'd0}, regs_4_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1546 = _T_1545 + _GEN_1760; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1761 = {{2'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1547 = _T_1546 + _GEN_1761; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1762 = {{3'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1548 = _T_1547 + _GEN_1762; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1763 = {{4'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1549 = _T_1548 + _GEN_1763; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1764 = {{5'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1550 = _T_1549 + _GEN_1764; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1765 = {{6'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1551 = _T_1550 + _GEN_1765; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1766 = {{7'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1552 = _T_1551 + _GEN_1766; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1767 = {{8'd0}, regs_5_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1554 = _T_1552 - _GEN_1767; // @[Conwaylife.scala 29:42]
  wire  _T_1555 = _T_1554 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1556 = _T_1554 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1557 = _T_1554 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1559 = regs_4_12 + regs_4_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1768 = {{1'd0}, regs_4_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1560 = _T_1559 + _GEN_1768; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1769 = {{2'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1561 = _T_1560 + _GEN_1769; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1770 = {{3'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1562 = _T_1561 + _GEN_1770; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1771 = {{4'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1563 = _T_1562 + _GEN_1771; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1772 = {{5'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1564 = _T_1563 + _GEN_1772; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1773 = {{6'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1565 = _T_1564 + _GEN_1773; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1774 = {{7'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1566 = _T_1565 + _GEN_1774; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1775 = {{8'd0}, regs_5_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1568 = _T_1566 - _GEN_1775; // @[Conwaylife.scala 29:42]
  wire  _T_1569 = _T_1568 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1570 = _T_1568 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1571 = _T_1568 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1573 = regs_4_13 + regs_4_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1776 = {{1'd0}, regs_4_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1574 = _T_1573 + _GEN_1776; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1777 = {{2'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1575 = _T_1574 + _GEN_1777; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1778 = {{3'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1576 = _T_1575 + _GEN_1778; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1779 = {{4'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1577 = _T_1576 + _GEN_1779; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1780 = {{5'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1578 = _T_1577 + _GEN_1780; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1781 = {{6'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1579 = _T_1578 + _GEN_1781; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1782 = {{7'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1580 = _T_1579 + _GEN_1782; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1783 = {{8'd0}, regs_5_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1582 = _T_1580 - _GEN_1783; // @[Conwaylife.scala 29:42]
  wire  _T_1583 = _T_1582 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1584 = _T_1582 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1585 = _T_1582 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1587 = regs_4_14 + regs_4_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1784 = {{1'd0}, regs_4_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1588 = _T_1587 + _GEN_1784; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1785 = {{2'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1589 = _T_1588 + _GEN_1785; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1786 = {{3'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1590 = _T_1589 + _GEN_1786; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1787 = {{4'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1591 = _T_1590 + _GEN_1787; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1788 = {{5'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1592 = _T_1591 + _GEN_1788; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1789 = {{6'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1593 = _T_1592 + _GEN_1789; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1790 = {{7'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1594 = _T_1593 + _GEN_1790; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1791 = {{8'd0}, regs_5_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1596 = _T_1594 - _GEN_1791; // @[Conwaylife.scala 29:42]
  wire  _T_1597 = _T_1596 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1598 = _T_1596 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1599 = _T_1596 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1601 = regs_5_15 + regs_5_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1792 = {{1'd0}, regs_5_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1602 = _T_1601 + _GEN_1792; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1793 = {{2'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1603 = _T_1602 + _GEN_1793; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1794 = {{3'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1604 = _T_1603 + _GEN_1794; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1795 = {{4'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1605 = _T_1604 + _GEN_1795; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1796 = {{5'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1606 = _T_1605 + _GEN_1796; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1797 = {{6'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1607 = _T_1606 + _GEN_1797; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1798 = {{7'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1608 = _T_1607 + _GEN_1798; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1799 = {{8'd0}, regs_6_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1610 = _T_1608 - _GEN_1799; // @[Conwaylife.scala 29:42]
  wire  _T_1611 = _T_1610 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1612 = _T_1610 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1613 = _T_1610 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1615 = regs_5_0 + regs_5_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1800 = {{1'd0}, regs_5_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1616 = _T_1615 + _GEN_1800; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1801 = {{2'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1617 = _T_1616 + _GEN_1801; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1802 = {{3'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1618 = _T_1617 + _GEN_1802; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1803 = {{4'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1619 = _T_1618 + _GEN_1803; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1804 = {{5'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1620 = _T_1619 + _GEN_1804; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1805 = {{6'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1621 = _T_1620 + _GEN_1805; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1806 = {{7'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1622 = _T_1621 + _GEN_1806; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1807 = {{8'd0}, regs_6_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1624 = _T_1622 - _GEN_1807; // @[Conwaylife.scala 29:42]
  wire  _T_1625 = _T_1624 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1626 = _T_1624 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1627 = _T_1624 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1629 = regs_5_1 + regs_5_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1808 = {{1'd0}, regs_5_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1630 = _T_1629 + _GEN_1808; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1809 = {{2'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1631 = _T_1630 + _GEN_1809; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1810 = {{3'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1632 = _T_1631 + _GEN_1810; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1811 = {{4'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1633 = _T_1632 + _GEN_1811; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1812 = {{5'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1634 = _T_1633 + _GEN_1812; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1813 = {{6'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1635 = _T_1634 + _GEN_1813; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1814 = {{7'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1636 = _T_1635 + _GEN_1814; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1815 = {{8'd0}, regs_6_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1638 = _T_1636 - _GEN_1815; // @[Conwaylife.scala 29:42]
  wire  _T_1639 = _T_1638 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1640 = _T_1638 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1641 = _T_1638 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1643 = regs_5_2 + regs_5_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1816 = {{1'd0}, regs_5_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1644 = _T_1643 + _GEN_1816; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1817 = {{2'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1645 = _T_1644 + _GEN_1817; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1818 = {{3'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1646 = _T_1645 + _GEN_1818; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1819 = {{4'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1647 = _T_1646 + _GEN_1819; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1820 = {{5'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1648 = _T_1647 + _GEN_1820; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1821 = {{6'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1649 = _T_1648 + _GEN_1821; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1822 = {{7'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1650 = _T_1649 + _GEN_1822; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1823 = {{8'd0}, regs_6_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1652 = _T_1650 - _GEN_1823; // @[Conwaylife.scala 29:42]
  wire  _T_1653 = _T_1652 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1654 = _T_1652 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1655 = _T_1652 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1657 = regs_5_3 + regs_5_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1824 = {{1'd0}, regs_5_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1658 = _T_1657 + _GEN_1824; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1825 = {{2'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1659 = _T_1658 + _GEN_1825; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1826 = {{3'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1660 = _T_1659 + _GEN_1826; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1827 = {{4'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1661 = _T_1660 + _GEN_1827; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1828 = {{5'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1662 = _T_1661 + _GEN_1828; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1829 = {{6'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1663 = _T_1662 + _GEN_1829; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1830 = {{7'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1664 = _T_1663 + _GEN_1830; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1831 = {{8'd0}, regs_6_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1666 = _T_1664 - _GEN_1831; // @[Conwaylife.scala 29:42]
  wire  _T_1667 = _T_1666 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1668 = _T_1666 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1669 = _T_1666 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1671 = regs_5_4 + regs_5_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1832 = {{1'd0}, regs_5_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1672 = _T_1671 + _GEN_1832; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1833 = {{2'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1673 = _T_1672 + _GEN_1833; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1834 = {{3'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1674 = _T_1673 + _GEN_1834; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1835 = {{4'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1675 = _T_1674 + _GEN_1835; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1836 = {{5'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1676 = _T_1675 + _GEN_1836; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1837 = {{6'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1677 = _T_1676 + _GEN_1837; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1838 = {{7'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1678 = _T_1677 + _GEN_1838; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1839 = {{8'd0}, regs_6_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1680 = _T_1678 - _GEN_1839; // @[Conwaylife.scala 29:42]
  wire  _T_1681 = _T_1680 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1682 = _T_1680 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1683 = _T_1680 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1685 = regs_5_5 + regs_5_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1840 = {{1'd0}, regs_5_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1686 = _T_1685 + _GEN_1840; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1841 = {{2'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1687 = _T_1686 + _GEN_1841; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1842 = {{3'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1688 = _T_1687 + _GEN_1842; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1843 = {{4'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1689 = _T_1688 + _GEN_1843; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1844 = {{5'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1690 = _T_1689 + _GEN_1844; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1845 = {{6'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1691 = _T_1690 + _GEN_1845; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1846 = {{7'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1692 = _T_1691 + _GEN_1846; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1847 = {{8'd0}, regs_6_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1694 = _T_1692 - _GEN_1847; // @[Conwaylife.scala 29:42]
  wire  _T_1695 = _T_1694 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1696 = _T_1694 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1697 = _T_1694 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1699 = regs_5_6 + regs_5_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1848 = {{1'd0}, regs_5_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1700 = _T_1699 + _GEN_1848; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1849 = {{2'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1701 = _T_1700 + _GEN_1849; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1850 = {{3'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1702 = _T_1701 + _GEN_1850; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1851 = {{4'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1703 = _T_1702 + _GEN_1851; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1852 = {{5'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1704 = _T_1703 + _GEN_1852; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1853 = {{6'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1705 = _T_1704 + _GEN_1853; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1854 = {{7'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1706 = _T_1705 + _GEN_1854; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1855 = {{8'd0}, regs_6_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1708 = _T_1706 - _GEN_1855; // @[Conwaylife.scala 29:42]
  wire  _T_1709 = _T_1708 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1710 = _T_1708 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1711 = _T_1708 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1713 = regs_5_7 + regs_5_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1856 = {{1'd0}, regs_5_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1714 = _T_1713 + _GEN_1856; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1857 = {{2'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1715 = _T_1714 + _GEN_1857; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1858 = {{3'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1716 = _T_1715 + _GEN_1858; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1859 = {{4'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1717 = _T_1716 + _GEN_1859; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1860 = {{5'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1718 = _T_1717 + _GEN_1860; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1861 = {{6'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1719 = _T_1718 + _GEN_1861; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1862 = {{7'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1720 = _T_1719 + _GEN_1862; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1863 = {{8'd0}, regs_6_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1722 = _T_1720 - _GEN_1863; // @[Conwaylife.scala 29:42]
  wire  _T_1723 = _T_1722 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1724 = _T_1722 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1725 = _T_1722 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1727 = regs_5_8 + regs_5_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1864 = {{1'd0}, regs_5_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1728 = _T_1727 + _GEN_1864; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1865 = {{2'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1729 = _T_1728 + _GEN_1865; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1866 = {{3'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1730 = _T_1729 + _GEN_1866; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1867 = {{4'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1731 = _T_1730 + _GEN_1867; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1868 = {{5'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1732 = _T_1731 + _GEN_1868; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1869 = {{6'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1733 = _T_1732 + _GEN_1869; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1870 = {{7'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1734 = _T_1733 + _GEN_1870; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1871 = {{8'd0}, regs_6_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1736 = _T_1734 - _GEN_1871; // @[Conwaylife.scala 29:42]
  wire  _T_1737 = _T_1736 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1738 = _T_1736 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1739 = _T_1736 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1741 = regs_5_9 + regs_5_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1872 = {{1'd0}, regs_5_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1742 = _T_1741 + _GEN_1872; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1873 = {{2'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1743 = _T_1742 + _GEN_1873; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1874 = {{3'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1744 = _T_1743 + _GEN_1874; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1875 = {{4'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1745 = _T_1744 + _GEN_1875; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1876 = {{5'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1746 = _T_1745 + _GEN_1876; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1877 = {{6'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1747 = _T_1746 + _GEN_1877; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1878 = {{7'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1748 = _T_1747 + _GEN_1878; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1879 = {{8'd0}, regs_6_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1750 = _T_1748 - _GEN_1879; // @[Conwaylife.scala 29:42]
  wire  _T_1751 = _T_1750 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1752 = _T_1750 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1753 = _T_1750 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1755 = regs_5_10 + regs_5_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1880 = {{1'd0}, regs_5_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1756 = _T_1755 + _GEN_1880; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1881 = {{2'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1757 = _T_1756 + _GEN_1881; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1882 = {{3'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1758 = _T_1757 + _GEN_1882; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1883 = {{4'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1759 = _T_1758 + _GEN_1883; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1884 = {{5'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1760 = _T_1759 + _GEN_1884; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1885 = {{6'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1761 = _T_1760 + _GEN_1885; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1886 = {{7'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1762 = _T_1761 + _GEN_1886; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1887 = {{8'd0}, regs_6_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1764 = _T_1762 - _GEN_1887; // @[Conwaylife.scala 29:42]
  wire  _T_1765 = _T_1764 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1766 = _T_1764 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1767 = _T_1764 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1769 = regs_5_11 + regs_5_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1888 = {{1'd0}, regs_5_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1770 = _T_1769 + _GEN_1888; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1889 = {{2'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1771 = _T_1770 + _GEN_1889; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1890 = {{3'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1772 = _T_1771 + _GEN_1890; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1891 = {{4'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1773 = _T_1772 + _GEN_1891; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1892 = {{5'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1774 = _T_1773 + _GEN_1892; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1893 = {{6'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1775 = _T_1774 + _GEN_1893; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1894 = {{7'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1776 = _T_1775 + _GEN_1894; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1895 = {{8'd0}, regs_6_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1778 = _T_1776 - _GEN_1895; // @[Conwaylife.scala 29:42]
  wire  _T_1779 = _T_1778 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1780 = _T_1778 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1781 = _T_1778 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1783 = regs_5_12 + regs_5_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1896 = {{1'd0}, regs_5_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1784 = _T_1783 + _GEN_1896; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1897 = {{2'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1785 = _T_1784 + _GEN_1897; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1898 = {{3'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1786 = _T_1785 + _GEN_1898; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1899 = {{4'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1787 = _T_1786 + _GEN_1899; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1900 = {{5'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1788 = _T_1787 + _GEN_1900; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1901 = {{6'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1789 = _T_1788 + _GEN_1901; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1902 = {{7'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1790 = _T_1789 + _GEN_1902; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1903 = {{8'd0}, regs_6_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1792 = _T_1790 - _GEN_1903; // @[Conwaylife.scala 29:42]
  wire  _T_1793 = _T_1792 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1794 = _T_1792 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1795 = _T_1792 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1797 = regs_5_13 + regs_5_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1904 = {{1'd0}, regs_5_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1798 = _T_1797 + _GEN_1904; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1905 = {{2'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1799 = _T_1798 + _GEN_1905; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1906 = {{3'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1800 = _T_1799 + _GEN_1906; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1907 = {{4'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1801 = _T_1800 + _GEN_1907; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1908 = {{5'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1802 = _T_1801 + _GEN_1908; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1909 = {{6'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1803 = _T_1802 + _GEN_1909; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1910 = {{7'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1804 = _T_1803 + _GEN_1910; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1911 = {{8'd0}, regs_6_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1806 = _T_1804 - _GEN_1911; // @[Conwaylife.scala 29:42]
  wire  _T_1807 = _T_1806 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1808 = _T_1806 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1809 = _T_1806 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1811 = regs_5_14 + regs_5_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1912 = {{1'd0}, regs_5_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1812 = _T_1811 + _GEN_1912; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1913 = {{2'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1813 = _T_1812 + _GEN_1913; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1914 = {{3'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1814 = _T_1813 + _GEN_1914; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1915 = {{4'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1815 = _T_1814 + _GEN_1915; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1916 = {{5'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1816 = _T_1815 + _GEN_1916; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1917 = {{6'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1817 = _T_1816 + _GEN_1917; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1918 = {{7'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1818 = _T_1817 + _GEN_1918; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1919 = {{8'd0}, regs_6_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1820 = _T_1818 - _GEN_1919; // @[Conwaylife.scala 29:42]
  wire  _T_1821 = _T_1820 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1822 = _T_1820 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1823 = _T_1820 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1825 = regs_6_15 + regs_6_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1920 = {{1'd0}, regs_6_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1826 = _T_1825 + _GEN_1920; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1921 = {{2'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1827 = _T_1826 + _GEN_1921; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1922 = {{3'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1828 = _T_1827 + _GEN_1922; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1923 = {{4'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1829 = _T_1828 + _GEN_1923; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1924 = {{5'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1830 = _T_1829 + _GEN_1924; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1925 = {{6'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1831 = _T_1830 + _GEN_1925; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1926 = {{7'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1832 = _T_1831 + _GEN_1926; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1927 = {{8'd0}, regs_7_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1834 = _T_1832 - _GEN_1927; // @[Conwaylife.scala 29:42]
  wire  _T_1835 = _T_1834 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1836 = _T_1834 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1837 = _T_1834 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1839 = regs_6_0 + regs_6_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1928 = {{1'd0}, regs_6_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1840 = _T_1839 + _GEN_1928; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1929 = {{2'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1841 = _T_1840 + _GEN_1929; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1930 = {{3'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1842 = _T_1841 + _GEN_1930; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1931 = {{4'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1843 = _T_1842 + _GEN_1931; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1932 = {{5'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1844 = _T_1843 + _GEN_1932; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1933 = {{6'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1845 = _T_1844 + _GEN_1933; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1934 = {{7'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1846 = _T_1845 + _GEN_1934; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1935 = {{8'd0}, regs_7_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1848 = _T_1846 - _GEN_1935; // @[Conwaylife.scala 29:42]
  wire  _T_1849 = _T_1848 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1850 = _T_1848 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1851 = _T_1848 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1853 = regs_6_1 + regs_6_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1936 = {{1'd0}, regs_6_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1854 = _T_1853 + _GEN_1936; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1937 = {{2'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1855 = _T_1854 + _GEN_1937; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1938 = {{3'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1856 = _T_1855 + _GEN_1938; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1939 = {{4'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1857 = _T_1856 + _GEN_1939; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1940 = {{5'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1858 = _T_1857 + _GEN_1940; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1941 = {{6'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1859 = _T_1858 + _GEN_1941; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1942 = {{7'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1860 = _T_1859 + _GEN_1942; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1943 = {{8'd0}, regs_7_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1862 = _T_1860 - _GEN_1943; // @[Conwaylife.scala 29:42]
  wire  _T_1863 = _T_1862 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1864 = _T_1862 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1865 = _T_1862 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1867 = regs_6_2 + regs_6_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1944 = {{1'd0}, regs_6_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1868 = _T_1867 + _GEN_1944; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1945 = {{2'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1869 = _T_1868 + _GEN_1945; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1946 = {{3'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1870 = _T_1869 + _GEN_1946; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1947 = {{4'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1871 = _T_1870 + _GEN_1947; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1948 = {{5'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1872 = _T_1871 + _GEN_1948; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1949 = {{6'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1873 = _T_1872 + _GEN_1949; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1950 = {{7'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1874 = _T_1873 + _GEN_1950; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1951 = {{8'd0}, regs_7_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1876 = _T_1874 - _GEN_1951; // @[Conwaylife.scala 29:42]
  wire  _T_1877 = _T_1876 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1878 = _T_1876 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1879 = _T_1876 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1881 = regs_6_3 + regs_6_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1952 = {{1'd0}, regs_6_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1882 = _T_1881 + _GEN_1952; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1953 = {{2'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1883 = _T_1882 + _GEN_1953; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1954 = {{3'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1884 = _T_1883 + _GEN_1954; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1955 = {{4'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1885 = _T_1884 + _GEN_1955; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1956 = {{5'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1886 = _T_1885 + _GEN_1956; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1957 = {{6'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1887 = _T_1886 + _GEN_1957; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1958 = {{7'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1888 = _T_1887 + _GEN_1958; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1959 = {{8'd0}, regs_7_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1890 = _T_1888 - _GEN_1959; // @[Conwaylife.scala 29:42]
  wire  _T_1891 = _T_1890 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1892 = _T_1890 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1893 = _T_1890 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1895 = regs_6_4 + regs_6_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1960 = {{1'd0}, regs_6_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1896 = _T_1895 + _GEN_1960; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1961 = {{2'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1897 = _T_1896 + _GEN_1961; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1962 = {{3'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1898 = _T_1897 + _GEN_1962; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1963 = {{4'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1899 = _T_1898 + _GEN_1963; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1964 = {{5'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1900 = _T_1899 + _GEN_1964; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1965 = {{6'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1901 = _T_1900 + _GEN_1965; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1966 = {{7'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1902 = _T_1901 + _GEN_1966; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1967 = {{8'd0}, regs_7_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1904 = _T_1902 - _GEN_1967; // @[Conwaylife.scala 29:42]
  wire  _T_1905 = _T_1904 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1906 = _T_1904 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1907 = _T_1904 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1909 = regs_6_5 + regs_6_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1968 = {{1'd0}, regs_6_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1910 = _T_1909 + _GEN_1968; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1969 = {{2'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1911 = _T_1910 + _GEN_1969; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1970 = {{3'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1912 = _T_1911 + _GEN_1970; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1971 = {{4'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1913 = _T_1912 + _GEN_1971; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1972 = {{5'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1914 = _T_1913 + _GEN_1972; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1973 = {{6'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1915 = _T_1914 + _GEN_1973; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1974 = {{7'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1916 = _T_1915 + _GEN_1974; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1975 = {{8'd0}, regs_7_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1918 = _T_1916 - _GEN_1975; // @[Conwaylife.scala 29:42]
  wire  _T_1919 = _T_1918 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1920 = _T_1918 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1921 = _T_1918 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1923 = regs_6_6 + regs_6_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1976 = {{1'd0}, regs_6_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1924 = _T_1923 + _GEN_1976; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1977 = {{2'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1925 = _T_1924 + _GEN_1977; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1978 = {{3'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1926 = _T_1925 + _GEN_1978; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1979 = {{4'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1927 = _T_1926 + _GEN_1979; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1980 = {{5'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1928 = _T_1927 + _GEN_1980; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1981 = {{6'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1929 = _T_1928 + _GEN_1981; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1982 = {{7'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1930 = _T_1929 + _GEN_1982; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1983 = {{8'd0}, regs_7_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1932 = _T_1930 - _GEN_1983; // @[Conwaylife.scala 29:42]
  wire  _T_1933 = _T_1932 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1934 = _T_1932 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1935 = _T_1932 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1937 = regs_6_7 + regs_6_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1984 = {{1'd0}, regs_6_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1938 = _T_1937 + _GEN_1984; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1985 = {{2'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1939 = _T_1938 + _GEN_1985; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1986 = {{3'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1940 = _T_1939 + _GEN_1986; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1987 = {{4'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1941 = _T_1940 + _GEN_1987; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1988 = {{5'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1942 = _T_1941 + _GEN_1988; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1989 = {{6'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1943 = _T_1942 + _GEN_1989; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1990 = {{7'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1944 = _T_1943 + _GEN_1990; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1991 = {{8'd0}, regs_7_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1946 = _T_1944 - _GEN_1991; // @[Conwaylife.scala 29:42]
  wire  _T_1947 = _T_1946 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1948 = _T_1946 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1949 = _T_1946 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1951 = regs_6_8 + regs_6_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_1992 = {{1'd0}, regs_6_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1952 = _T_1951 + _GEN_1992; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_1993 = {{2'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1953 = _T_1952 + _GEN_1993; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_1994 = {{3'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1954 = _T_1953 + _GEN_1994; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_1995 = {{4'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1955 = _T_1954 + _GEN_1995; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_1996 = {{5'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1956 = _T_1955 + _GEN_1996; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_1997 = {{6'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1957 = _T_1956 + _GEN_1997; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_1998 = {{7'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1958 = _T_1957 + _GEN_1998; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_1999 = {{8'd0}, regs_7_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1960 = _T_1958 - _GEN_1999; // @[Conwaylife.scala 29:42]
  wire  _T_1961 = _T_1960 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1962 = _T_1960 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1963 = _T_1960 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1965 = regs_6_9 + regs_6_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2000 = {{1'd0}, regs_6_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1966 = _T_1965 + _GEN_2000; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2001 = {{2'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1967 = _T_1966 + _GEN_2001; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2002 = {{3'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1968 = _T_1967 + _GEN_2002; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2003 = {{4'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1969 = _T_1968 + _GEN_2003; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2004 = {{5'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1970 = _T_1969 + _GEN_2004; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2005 = {{6'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1971 = _T_1970 + _GEN_2005; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2006 = {{7'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1972 = _T_1971 + _GEN_2006; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2007 = {{8'd0}, regs_7_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1974 = _T_1972 - _GEN_2007; // @[Conwaylife.scala 29:42]
  wire  _T_1975 = _T_1974 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1976 = _T_1974 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1977 = _T_1974 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1979 = regs_6_10 + regs_6_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2008 = {{1'd0}, regs_6_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1980 = _T_1979 + _GEN_2008; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2009 = {{2'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1981 = _T_1980 + _GEN_2009; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2010 = {{3'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1982 = _T_1981 + _GEN_2010; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2011 = {{4'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1983 = _T_1982 + _GEN_2011; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2012 = {{5'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1984 = _T_1983 + _GEN_2012; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2013 = {{6'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1985 = _T_1984 + _GEN_2013; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2014 = {{7'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_1986 = _T_1985 + _GEN_2014; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2015 = {{8'd0}, regs_7_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_1988 = _T_1986 - _GEN_2015; // @[Conwaylife.scala 29:42]
  wire  _T_1989 = _T_1988 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_1990 = _T_1988 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_1991 = _T_1988 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_1993 = regs_6_11 + regs_6_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2016 = {{1'd0}, regs_6_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_1994 = _T_1993 + _GEN_2016; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2017 = {{2'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_1995 = _T_1994 + _GEN_2017; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2018 = {{3'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_1996 = _T_1995 + _GEN_2018; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2019 = {{4'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_1997 = _T_1996 + _GEN_2019; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2020 = {{5'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_1998 = _T_1997 + _GEN_2020; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2021 = {{6'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_1999 = _T_1998 + _GEN_2021; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2022 = {{7'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2000 = _T_1999 + _GEN_2022; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2023 = {{8'd0}, regs_7_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2002 = _T_2000 - _GEN_2023; // @[Conwaylife.scala 29:42]
  wire  _T_2003 = _T_2002 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2004 = _T_2002 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2005 = _T_2002 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2007 = regs_6_12 + regs_6_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2024 = {{1'd0}, regs_6_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2008 = _T_2007 + _GEN_2024; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2025 = {{2'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2009 = _T_2008 + _GEN_2025; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2026 = {{3'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2010 = _T_2009 + _GEN_2026; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2027 = {{4'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2011 = _T_2010 + _GEN_2027; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2028 = {{5'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2012 = _T_2011 + _GEN_2028; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2029 = {{6'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2013 = _T_2012 + _GEN_2029; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2030 = {{7'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2014 = _T_2013 + _GEN_2030; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2031 = {{8'd0}, regs_7_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2016 = _T_2014 - _GEN_2031; // @[Conwaylife.scala 29:42]
  wire  _T_2017 = _T_2016 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2018 = _T_2016 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2019 = _T_2016 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2021 = regs_6_13 + regs_6_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2032 = {{1'd0}, regs_6_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2022 = _T_2021 + _GEN_2032; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2033 = {{2'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2023 = _T_2022 + _GEN_2033; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2034 = {{3'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2024 = _T_2023 + _GEN_2034; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2035 = {{4'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2025 = _T_2024 + _GEN_2035; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2036 = {{5'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2026 = _T_2025 + _GEN_2036; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2037 = {{6'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2027 = _T_2026 + _GEN_2037; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2038 = {{7'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2028 = _T_2027 + _GEN_2038; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2039 = {{8'd0}, regs_7_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2030 = _T_2028 - _GEN_2039; // @[Conwaylife.scala 29:42]
  wire  _T_2031 = _T_2030 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2032 = _T_2030 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2033 = _T_2030 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2035 = regs_6_14 + regs_6_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2040 = {{1'd0}, regs_6_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2036 = _T_2035 + _GEN_2040; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2041 = {{2'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2037 = _T_2036 + _GEN_2041; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2042 = {{3'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2038 = _T_2037 + _GEN_2042; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2043 = {{4'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2039 = _T_2038 + _GEN_2043; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2044 = {{5'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2040 = _T_2039 + _GEN_2044; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2045 = {{6'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2041 = _T_2040 + _GEN_2045; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2046 = {{7'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2042 = _T_2041 + _GEN_2046; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2047 = {{8'd0}, regs_7_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2044 = _T_2042 - _GEN_2047; // @[Conwaylife.scala 29:42]
  wire  _T_2045 = _T_2044 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2046 = _T_2044 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2047 = _T_2044 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2049 = regs_7_15 + regs_7_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2048 = {{1'd0}, regs_7_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2050 = _T_2049 + _GEN_2048; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2049 = {{2'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2051 = _T_2050 + _GEN_2049; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2050 = {{3'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2052 = _T_2051 + _GEN_2050; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2051 = {{4'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2053 = _T_2052 + _GEN_2051; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2052 = {{5'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2054 = _T_2053 + _GEN_2052; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2053 = {{6'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2055 = _T_2054 + _GEN_2053; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2054 = {{7'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2056 = _T_2055 + _GEN_2054; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2055 = {{8'd0}, regs_8_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2058 = _T_2056 - _GEN_2055; // @[Conwaylife.scala 29:42]
  wire  _T_2059 = _T_2058 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2060 = _T_2058 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2061 = _T_2058 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2063 = regs_7_0 + regs_7_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2056 = {{1'd0}, regs_7_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2064 = _T_2063 + _GEN_2056; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2057 = {{2'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2065 = _T_2064 + _GEN_2057; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2058 = {{3'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2066 = _T_2065 + _GEN_2058; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2059 = {{4'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2067 = _T_2066 + _GEN_2059; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2060 = {{5'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2068 = _T_2067 + _GEN_2060; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2061 = {{6'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2069 = _T_2068 + _GEN_2061; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2062 = {{7'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2070 = _T_2069 + _GEN_2062; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2063 = {{8'd0}, regs_8_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2072 = _T_2070 - _GEN_2063; // @[Conwaylife.scala 29:42]
  wire  _T_2073 = _T_2072 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2074 = _T_2072 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2075 = _T_2072 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2077 = regs_7_1 + regs_7_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2064 = {{1'd0}, regs_7_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2078 = _T_2077 + _GEN_2064; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2065 = {{2'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2079 = _T_2078 + _GEN_2065; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2066 = {{3'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2080 = _T_2079 + _GEN_2066; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2067 = {{4'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2081 = _T_2080 + _GEN_2067; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2068 = {{5'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2082 = _T_2081 + _GEN_2068; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2069 = {{6'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2083 = _T_2082 + _GEN_2069; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2070 = {{7'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2084 = _T_2083 + _GEN_2070; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2071 = {{8'd0}, regs_8_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2086 = _T_2084 - _GEN_2071; // @[Conwaylife.scala 29:42]
  wire  _T_2087 = _T_2086 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2088 = _T_2086 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2089 = _T_2086 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2091 = regs_7_2 + regs_7_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2072 = {{1'd0}, regs_7_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2092 = _T_2091 + _GEN_2072; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2073 = {{2'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2093 = _T_2092 + _GEN_2073; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2074 = {{3'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2094 = _T_2093 + _GEN_2074; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2075 = {{4'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2095 = _T_2094 + _GEN_2075; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2076 = {{5'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2096 = _T_2095 + _GEN_2076; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2077 = {{6'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2097 = _T_2096 + _GEN_2077; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2078 = {{7'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2098 = _T_2097 + _GEN_2078; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2079 = {{8'd0}, regs_8_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2100 = _T_2098 - _GEN_2079; // @[Conwaylife.scala 29:42]
  wire  _T_2101 = _T_2100 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2102 = _T_2100 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2103 = _T_2100 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2105 = regs_7_3 + regs_7_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2080 = {{1'd0}, regs_7_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2106 = _T_2105 + _GEN_2080; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2081 = {{2'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2107 = _T_2106 + _GEN_2081; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2082 = {{3'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2108 = _T_2107 + _GEN_2082; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2083 = {{4'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2109 = _T_2108 + _GEN_2083; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2084 = {{5'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2110 = _T_2109 + _GEN_2084; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2085 = {{6'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2111 = _T_2110 + _GEN_2085; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2086 = {{7'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2112 = _T_2111 + _GEN_2086; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2087 = {{8'd0}, regs_8_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2114 = _T_2112 - _GEN_2087; // @[Conwaylife.scala 29:42]
  wire  _T_2115 = _T_2114 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2116 = _T_2114 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2117 = _T_2114 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2119 = regs_7_4 + regs_7_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2088 = {{1'd0}, regs_7_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2120 = _T_2119 + _GEN_2088; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2089 = {{2'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2121 = _T_2120 + _GEN_2089; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2090 = {{3'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2122 = _T_2121 + _GEN_2090; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2091 = {{4'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2123 = _T_2122 + _GEN_2091; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2092 = {{5'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2124 = _T_2123 + _GEN_2092; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2093 = {{6'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2125 = _T_2124 + _GEN_2093; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2094 = {{7'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2126 = _T_2125 + _GEN_2094; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2095 = {{8'd0}, regs_8_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2128 = _T_2126 - _GEN_2095; // @[Conwaylife.scala 29:42]
  wire  _T_2129 = _T_2128 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2130 = _T_2128 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2131 = _T_2128 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2133 = regs_7_5 + regs_7_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2096 = {{1'd0}, regs_7_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2134 = _T_2133 + _GEN_2096; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2097 = {{2'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2135 = _T_2134 + _GEN_2097; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2098 = {{3'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2136 = _T_2135 + _GEN_2098; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2099 = {{4'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2137 = _T_2136 + _GEN_2099; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2100 = {{5'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2138 = _T_2137 + _GEN_2100; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2101 = {{6'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2139 = _T_2138 + _GEN_2101; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2102 = {{7'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2140 = _T_2139 + _GEN_2102; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2103 = {{8'd0}, regs_8_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2142 = _T_2140 - _GEN_2103; // @[Conwaylife.scala 29:42]
  wire  _T_2143 = _T_2142 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2144 = _T_2142 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2145 = _T_2142 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2147 = regs_7_6 + regs_7_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2104 = {{1'd0}, regs_7_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2148 = _T_2147 + _GEN_2104; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2105 = {{2'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2149 = _T_2148 + _GEN_2105; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2106 = {{3'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2150 = _T_2149 + _GEN_2106; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2107 = {{4'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2151 = _T_2150 + _GEN_2107; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2108 = {{5'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2152 = _T_2151 + _GEN_2108; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2109 = {{6'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2153 = _T_2152 + _GEN_2109; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2110 = {{7'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2154 = _T_2153 + _GEN_2110; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2111 = {{8'd0}, regs_8_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2156 = _T_2154 - _GEN_2111; // @[Conwaylife.scala 29:42]
  wire  _T_2157 = _T_2156 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2158 = _T_2156 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2159 = _T_2156 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2161 = regs_7_7 + regs_7_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2112 = {{1'd0}, regs_7_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2162 = _T_2161 + _GEN_2112; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2113 = {{2'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2163 = _T_2162 + _GEN_2113; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2114 = {{3'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2164 = _T_2163 + _GEN_2114; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2115 = {{4'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2165 = _T_2164 + _GEN_2115; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2116 = {{5'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2166 = _T_2165 + _GEN_2116; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2117 = {{6'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2167 = _T_2166 + _GEN_2117; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2118 = {{7'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2168 = _T_2167 + _GEN_2118; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2119 = {{8'd0}, regs_8_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2170 = _T_2168 - _GEN_2119; // @[Conwaylife.scala 29:42]
  wire  _T_2171 = _T_2170 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2172 = _T_2170 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2173 = _T_2170 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2175 = regs_7_8 + regs_7_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2120 = {{1'd0}, regs_7_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2176 = _T_2175 + _GEN_2120; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2121 = {{2'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2177 = _T_2176 + _GEN_2121; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2122 = {{3'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2178 = _T_2177 + _GEN_2122; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2123 = {{4'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2179 = _T_2178 + _GEN_2123; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2124 = {{5'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2180 = _T_2179 + _GEN_2124; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2125 = {{6'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2181 = _T_2180 + _GEN_2125; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2126 = {{7'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2182 = _T_2181 + _GEN_2126; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2127 = {{8'd0}, regs_8_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2184 = _T_2182 - _GEN_2127; // @[Conwaylife.scala 29:42]
  wire  _T_2185 = _T_2184 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2186 = _T_2184 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2187 = _T_2184 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2189 = regs_7_9 + regs_7_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2128 = {{1'd0}, regs_7_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2190 = _T_2189 + _GEN_2128; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2129 = {{2'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2191 = _T_2190 + _GEN_2129; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2130 = {{3'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2192 = _T_2191 + _GEN_2130; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2131 = {{4'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2193 = _T_2192 + _GEN_2131; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2132 = {{5'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2194 = _T_2193 + _GEN_2132; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2133 = {{6'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2195 = _T_2194 + _GEN_2133; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2134 = {{7'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2196 = _T_2195 + _GEN_2134; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2135 = {{8'd0}, regs_8_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2198 = _T_2196 - _GEN_2135; // @[Conwaylife.scala 29:42]
  wire  _T_2199 = _T_2198 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2200 = _T_2198 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2201 = _T_2198 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2203 = regs_7_10 + regs_7_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2136 = {{1'd0}, regs_7_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2204 = _T_2203 + _GEN_2136; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2137 = {{2'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2205 = _T_2204 + _GEN_2137; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2138 = {{3'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2206 = _T_2205 + _GEN_2138; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2139 = {{4'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2207 = _T_2206 + _GEN_2139; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2140 = {{5'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2208 = _T_2207 + _GEN_2140; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2141 = {{6'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2209 = _T_2208 + _GEN_2141; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2142 = {{7'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2210 = _T_2209 + _GEN_2142; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2143 = {{8'd0}, regs_8_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2212 = _T_2210 - _GEN_2143; // @[Conwaylife.scala 29:42]
  wire  _T_2213 = _T_2212 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2214 = _T_2212 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2215 = _T_2212 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2217 = regs_7_11 + regs_7_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2144 = {{1'd0}, regs_7_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2218 = _T_2217 + _GEN_2144; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2145 = {{2'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2219 = _T_2218 + _GEN_2145; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2146 = {{3'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2220 = _T_2219 + _GEN_2146; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2147 = {{4'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2221 = _T_2220 + _GEN_2147; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2148 = {{5'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2222 = _T_2221 + _GEN_2148; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2149 = {{6'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2223 = _T_2222 + _GEN_2149; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2150 = {{7'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2224 = _T_2223 + _GEN_2150; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2151 = {{8'd0}, regs_8_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2226 = _T_2224 - _GEN_2151; // @[Conwaylife.scala 29:42]
  wire  _T_2227 = _T_2226 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2228 = _T_2226 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2229 = _T_2226 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2231 = regs_7_12 + regs_7_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2152 = {{1'd0}, regs_7_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2232 = _T_2231 + _GEN_2152; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2153 = {{2'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2233 = _T_2232 + _GEN_2153; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2154 = {{3'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2234 = _T_2233 + _GEN_2154; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2155 = {{4'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2235 = _T_2234 + _GEN_2155; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2156 = {{5'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2236 = _T_2235 + _GEN_2156; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2157 = {{6'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2237 = _T_2236 + _GEN_2157; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2158 = {{7'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2238 = _T_2237 + _GEN_2158; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2159 = {{8'd0}, regs_8_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2240 = _T_2238 - _GEN_2159; // @[Conwaylife.scala 29:42]
  wire  _T_2241 = _T_2240 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2242 = _T_2240 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2243 = _T_2240 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2245 = regs_7_13 + regs_7_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2160 = {{1'd0}, regs_7_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2246 = _T_2245 + _GEN_2160; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2161 = {{2'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2247 = _T_2246 + _GEN_2161; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2162 = {{3'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2248 = _T_2247 + _GEN_2162; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2163 = {{4'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2249 = _T_2248 + _GEN_2163; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2164 = {{5'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2250 = _T_2249 + _GEN_2164; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2165 = {{6'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2251 = _T_2250 + _GEN_2165; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2166 = {{7'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2252 = _T_2251 + _GEN_2166; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2167 = {{8'd0}, regs_8_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2254 = _T_2252 - _GEN_2167; // @[Conwaylife.scala 29:42]
  wire  _T_2255 = _T_2254 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2256 = _T_2254 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2257 = _T_2254 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2259 = regs_7_14 + regs_7_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2168 = {{1'd0}, regs_7_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2260 = _T_2259 + _GEN_2168; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2169 = {{2'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2261 = _T_2260 + _GEN_2169; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2170 = {{3'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2262 = _T_2261 + _GEN_2170; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2171 = {{4'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2263 = _T_2262 + _GEN_2171; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2172 = {{5'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2264 = _T_2263 + _GEN_2172; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2173 = {{6'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2265 = _T_2264 + _GEN_2173; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2174 = {{7'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2266 = _T_2265 + _GEN_2174; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2175 = {{8'd0}, regs_8_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2268 = _T_2266 - _GEN_2175; // @[Conwaylife.scala 29:42]
  wire  _T_2269 = _T_2268 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2270 = _T_2268 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2271 = _T_2268 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2273 = regs_8_15 + regs_8_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2176 = {{1'd0}, regs_8_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2274 = _T_2273 + _GEN_2176; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2177 = {{2'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2275 = _T_2274 + _GEN_2177; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2178 = {{3'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2276 = _T_2275 + _GEN_2178; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2179 = {{4'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2277 = _T_2276 + _GEN_2179; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2180 = {{5'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2278 = _T_2277 + _GEN_2180; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2181 = {{6'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2279 = _T_2278 + _GEN_2181; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2182 = {{7'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2280 = _T_2279 + _GEN_2182; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2183 = {{8'd0}, regs_9_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2282 = _T_2280 - _GEN_2183; // @[Conwaylife.scala 29:42]
  wire  _T_2283 = _T_2282 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2284 = _T_2282 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2285 = _T_2282 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2287 = regs_8_0 + regs_8_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2184 = {{1'd0}, regs_8_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2288 = _T_2287 + _GEN_2184; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2185 = {{2'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2289 = _T_2288 + _GEN_2185; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2186 = {{3'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2290 = _T_2289 + _GEN_2186; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2187 = {{4'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2291 = _T_2290 + _GEN_2187; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2188 = {{5'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2292 = _T_2291 + _GEN_2188; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2189 = {{6'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2293 = _T_2292 + _GEN_2189; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2190 = {{7'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2294 = _T_2293 + _GEN_2190; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2191 = {{8'd0}, regs_9_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2296 = _T_2294 - _GEN_2191; // @[Conwaylife.scala 29:42]
  wire  _T_2297 = _T_2296 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2298 = _T_2296 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2299 = _T_2296 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2301 = regs_8_1 + regs_8_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2192 = {{1'd0}, regs_8_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2302 = _T_2301 + _GEN_2192; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2193 = {{2'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2303 = _T_2302 + _GEN_2193; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2194 = {{3'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2304 = _T_2303 + _GEN_2194; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2195 = {{4'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2305 = _T_2304 + _GEN_2195; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2196 = {{5'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2306 = _T_2305 + _GEN_2196; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2197 = {{6'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2307 = _T_2306 + _GEN_2197; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2198 = {{7'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2308 = _T_2307 + _GEN_2198; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2199 = {{8'd0}, regs_9_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2310 = _T_2308 - _GEN_2199; // @[Conwaylife.scala 29:42]
  wire  _T_2311 = _T_2310 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2312 = _T_2310 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2313 = _T_2310 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2315 = regs_8_2 + regs_8_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2200 = {{1'd0}, regs_8_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2316 = _T_2315 + _GEN_2200; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2201 = {{2'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2317 = _T_2316 + _GEN_2201; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2202 = {{3'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2318 = _T_2317 + _GEN_2202; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2203 = {{4'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2319 = _T_2318 + _GEN_2203; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2204 = {{5'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2320 = _T_2319 + _GEN_2204; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2205 = {{6'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2321 = _T_2320 + _GEN_2205; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2206 = {{7'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2322 = _T_2321 + _GEN_2206; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2207 = {{8'd0}, regs_9_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2324 = _T_2322 - _GEN_2207; // @[Conwaylife.scala 29:42]
  wire  _T_2325 = _T_2324 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2326 = _T_2324 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2327 = _T_2324 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2329 = regs_8_3 + regs_8_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2208 = {{1'd0}, regs_8_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2330 = _T_2329 + _GEN_2208; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2209 = {{2'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2331 = _T_2330 + _GEN_2209; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2210 = {{3'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2332 = _T_2331 + _GEN_2210; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2211 = {{4'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2333 = _T_2332 + _GEN_2211; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2212 = {{5'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2334 = _T_2333 + _GEN_2212; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2213 = {{6'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2335 = _T_2334 + _GEN_2213; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2214 = {{7'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2336 = _T_2335 + _GEN_2214; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2215 = {{8'd0}, regs_9_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2338 = _T_2336 - _GEN_2215; // @[Conwaylife.scala 29:42]
  wire  _T_2339 = _T_2338 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2340 = _T_2338 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2341 = _T_2338 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2343 = regs_8_4 + regs_8_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2216 = {{1'd0}, regs_8_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2344 = _T_2343 + _GEN_2216; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2217 = {{2'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2345 = _T_2344 + _GEN_2217; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2218 = {{3'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2346 = _T_2345 + _GEN_2218; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2219 = {{4'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2347 = _T_2346 + _GEN_2219; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2220 = {{5'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2348 = _T_2347 + _GEN_2220; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2221 = {{6'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2349 = _T_2348 + _GEN_2221; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2222 = {{7'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2350 = _T_2349 + _GEN_2222; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2223 = {{8'd0}, regs_9_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2352 = _T_2350 - _GEN_2223; // @[Conwaylife.scala 29:42]
  wire  _T_2353 = _T_2352 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2354 = _T_2352 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2355 = _T_2352 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2357 = regs_8_5 + regs_8_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2224 = {{1'd0}, regs_8_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2358 = _T_2357 + _GEN_2224; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2225 = {{2'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2359 = _T_2358 + _GEN_2225; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2226 = {{3'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2360 = _T_2359 + _GEN_2226; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2227 = {{4'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2361 = _T_2360 + _GEN_2227; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2228 = {{5'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2362 = _T_2361 + _GEN_2228; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2229 = {{6'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2363 = _T_2362 + _GEN_2229; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2230 = {{7'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2364 = _T_2363 + _GEN_2230; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2231 = {{8'd0}, regs_9_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2366 = _T_2364 - _GEN_2231; // @[Conwaylife.scala 29:42]
  wire  _T_2367 = _T_2366 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2368 = _T_2366 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2369 = _T_2366 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2371 = regs_8_6 + regs_8_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2232 = {{1'd0}, regs_8_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2372 = _T_2371 + _GEN_2232; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2233 = {{2'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2373 = _T_2372 + _GEN_2233; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2234 = {{3'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2374 = _T_2373 + _GEN_2234; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2235 = {{4'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2375 = _T_2374 + _GEN_2235; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2236 = {{5'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2376 = _T_2375 + _GEN_2236; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2237 = {{6'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2377 = _T_2376 + _GEN_2237; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2238 = {{7'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2378 = _T_2377 + _GEN_2238; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2239 = {{8'd0}, regs_9_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2380 = _T_2378 - _GEN_2239; // @[Conwaylife.scala 29:42]
  wire  _T_2381 = _T_2380 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2382 = _T_2380 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2383 = _T_2380 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2385 = regs_8_7 + regs_8_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2240 = {{1'd0}, regs_8_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2386 = _T_2385 + _GEN_2240; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2241 = {{2'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2387 = _T_2386 + _GEN_2241; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2242 = {{3'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2388 = _T_2387 + _GEN_2242; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2243 = {{4'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2389 = _T_2388 + _GEN_2243; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2244 = {{5'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2390 = _T_2389 + _GEN_2244; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2245 = {{6'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2391 = _T_2390 + _GEN_2245; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2246 = {{7'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2392 = _T_2391 + _GEN_2246; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2247 = {{8'd0}, regs_9_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2394 = _T_2392 - _GEN_2247; // @[Conwaylife.scala 29:42]
  wire  _T_2395 = _T_2394 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2396 = _T_2394 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2397 = _T_2394 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2399 = regs_8_8 + regs_8_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2248 = {{1'd0}, regs_8_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2400 = _T_2399 + _GEN_2248; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2249 = {{2'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2401 = _T_2400 + _GEN_2249; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2250 = {{3'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2402 = _T_2401 + _GEN_2250; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2251 = {{4'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2403 = _T_2402 + _GEN_2251; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2252 = {{5'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2404 = _T_2403 + _GEN_2252; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2253 = {{6'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2405 = _T_2404 + _GEN_2253; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2254 = {{7'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2406 = _T_2405 + _GEN_2254; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2255 = {{8'd0}, regs_9_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2408 = _T_2406 - _GEN_2255; // @[Conwaylife.scala 29:42]
  wire  _T_2409 = _T_2408 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2410 = _T_2408 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2411 = _T_2408 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2413 = regs_8_9 + regs_8_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2256 = {{1'd0}, regs_8_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2414 = _T_2413 + _GEN_2256; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2257 = {{2'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2415 = _T_2414 + _GEN_2257; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2258 = {{3'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2416 = _T_2415 + _GEN_2258; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2259 = {{4'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2417 = _T_2416 + _GEN_2259; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2260 = {{5'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2418 = _T_2417 + _GEN_2260; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2261 = {{6'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2419 = _T_2418 + _GEN_2261; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2262 = {{7'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2420 = _T_2419 + _GEN_2262; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2263 = {{8'd0}, regs_9_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2422 = _T_2420 - _GEN_2263; // @[Conwaylife.scala 29:42]
  wire  _T_2423 = _T_2422 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2424 = _T_2422 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2425 = _T_2422 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2427 = regs_8_10 + regs_8_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2264 = {{1'd0}, regs_8_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2428 = _T_2427 + _GEN_2264; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2265 = {{2'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2429 = _T_2428 + _GEN_2265; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2266 = {{3'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2430 = _T_2429 + _GEN_2266; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2267 = {{4'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2431 = _T_2430 + _GEN_2267; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2268 = {{5'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2432 = _T_2431 + _GEN_2268; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2269 = {{6'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2433 = _T_2432 + _GEN_2269; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2270 = {{7'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2434 = _T_2433 + _GEN_2270; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2271 = {{8'd0}, regs_9_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2436 = _T_2434 - _GEN_2271; // @[Conwaylife.scala 29:42]
  wire  _T_2437 = _T_2436 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2438 = _T_2436 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2439 = _T_2436 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2441 = regs_8_11 + regs_8_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2272 = {{1'd0}, regs_8_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2442 = _T_2441 + _GEN_2272; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2273 = {{2'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2443 = _T_2442 + _GEN_2273; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2274 = {{3'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2444 = _T_2443 + _GEN_2274; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2275 = {{4'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2445 = _T_2444 + _GEN_2275; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2276 = {{5'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2446 = _T_2445 + _GEN_2276; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2277 = {{6'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2447 = _T_2446 + _GEN_2277; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2278 = {{7'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2448 = _T_2447 + _GEN_2278; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2279 = {{8'd0}, regs_9_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2450 = _T_2448 - _GEN_2279; // @[Conwaylife.scala 29:42]
  wire  _T_2451 = _T_2450 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2452 = _T_2450 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2453 = _T_2450 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2455 = regs_8_12 + regs_8_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2280 = {{1'd0}, regs_8_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2456 = _T_2455 + _GEN_2280; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2281 = {{2'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2457 = _T_2456 + _GEN_2281; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2282 = {{3'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2458 = _T_2457 + _GEN_2282; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2283 = {{4'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2459 = _T_2458 + _GEN_2283; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2284 = {{5'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2460 = _T_2459 + _GEN_2284; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2285 = {{6'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2461 = _T_2460 + _GEN_2285; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2286 = {{7'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2462 = _T_2461 + _GEN_2286; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2287 = {{8'd0}, regs_9_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2464 = _T_2462 - _GEN_2287; // @[Conwaylife.scala 29:42]
  wire  _T_2465 = _T_2464 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2466 = _T_2464 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2467 = _T_2464 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2469 = regs_8_13 + regs_8_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2288 = {{1'd0}, regs_8_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2470 = _T_2469 + _GEN_2288; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2289 = {{2'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2471 = _T_2470 + _GEN_2289; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2290 = {{3'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2472 = _T_2471 + _GEN_2290; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2291 = {{4'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2473 = _T_2472 + _GEN_2291; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2292 = {{5'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2474 = _T_2473 + _GEN_2292; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2293 = {{6'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2475 = _T_2474 + _GEN_2293; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2294 = {{7'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2476 = _T_2475 + _GEN_2294; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2295 = {{8'd0}, regs_9_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2478 = _T_2476 - _GEN_2295; // @[Conwaylife.scala 29:42]
  wire  _T_2479 = _T_2478 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2480 = _T_2478 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2481 = _T_2478 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2483 = regs_8_14 + regs_8_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2296 = {{1'd0}, regs_8_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2484 = _T_2483 + _GEN_2296; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2297 = {{2'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2485 = _T_2484 + _GEN_2297; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2298 = {{3'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2486 = _T_2485 + _GEN_2298; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2299 = {{4'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2487 = _T_2486 + _GEN_2299; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2300 = {{5'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2488 = _T_2487 + _GEN_2300; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2301 = {{6'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2489 = _T_2488 + _GEN_2301; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2302 = {{7'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2490 = _T_2489 + _GEN_2302; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2303 = {{8'd0}, regs_9_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2492 = _T_2490 - _GEN_2303; // @[Conwaylife.scala 29:42]
  wire  _T_2493 = _T_2492 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2494 = _T_2492 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2495 = _T_2492 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2497 = regs_9_15 + regs_9_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2304 = {{1'd0}, regs_9_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2498 = _T_2497 + _GEN_2304; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2305 = {{2'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2499 = _T_2498 + _GEN_2305; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2306 = {{3'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2500 = _T_2499 + _GEN_2306; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2307 = {{4'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2501 = _T_2500 + _GEN_2307; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2308 = {{5'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2502 = _T_2501 + _GEN_2308; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2309 = {{6'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2503 = _T_2502 + _GEN_2309; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2310 = {{7'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2504 = _T_2503 + _GEN_2310; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2311 = {{8'd0}, regs_10_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2506 = _T_2504 - _GEN_2311; // @[Conwaylife.scala 29:42]
  wire  _T_2507 = _T_2506 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2508 = _T_2506 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2509 = _T_2506 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2511 = regs_9_0 + regs_9_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2312 = {{1'd0}, regs_9_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2512 = _T_2511 + _GEN_2312; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2313 = {{2'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2513 = _T_2512 + _GEN_2313; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2314 = {{3'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2514 = _T_2513 + _GEN_2314; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2315 = {{4'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2515 = _T_2514 + _GEN_2315; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2316 = {{5'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2516 = _T_2515 + _GEN_2316; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2317 = {{6'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2517 = _T_2516 + _GEN_2317; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2318 = {{7'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2518 = _T_2517 + _GEN_2318; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2319 = {{8'd0}, regs_10_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2520 = _T_2518 - _GEN_2319; // @[Conwaylife.scala 29:42]
  wire  _T_2521 = _T_2520 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2522 = _T_2520 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2523 = _T_2520 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2525 = regs_9_1 + regs_9_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2320 = {{1'd0}, regs_9_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2526 = _T_2525 + _GEN_2320; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2321 = {{2'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2527 = _T_2526 + _GEN_2321; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2322 = {{3'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2528 = _T_2527 + _GEN_2322; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2323 = {{4'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2529 = _T_2528 + _GEN_2323; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2324 = {{5'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2530 = _T_2529 + _GEN_2324; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2325 = {{6'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2531 = _T_2530 + _GEN_2325; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2326 = {{7'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2532 = _T_2531 + _GEN_2326; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2327 = {{8'd0}, regs_10_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2534 = _T_2532 - _GEN_2327; // @[Conwaylife.scala 29:42]
  wire  _T_2535 = _T_2534 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2536 = _T_2534 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2537 = _T_2534 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2539 = regs_9_2 + regs_9_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2328 = {{1'd0}, regs_9_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2540 = _T_2539 + _GEN_2328; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2329 = {{2'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2541 = _T_2540 + _GEN_2329; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2330 = {{3'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2542 = _T_2541 + _GEN_2330; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2331 = {{4'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2543 = _T_2542 + _GEN_2331; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2332 = {{5'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2544 = _T_2543 + _GEN_2332; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2333 = {{6'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2545 = _T_2544 + _GEN_2333; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2334 = {{7'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2546 = _T_2545 + _GEN_2334; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2335 = {{8'd0}, regs_10_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2548 = _T_2546 - _GEN_2335; // @[Conwaylife.scala 29:42]
  wire  _T_2549 = _T_2548 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2550 = _T_2548 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2551 = _T_2548 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2553 = regs_9_3 + regs_9_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2336 = {{1'd0}, regs_9_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2554 = _T_2553 + _GEN_2336; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2337 = {{2'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2555 = _T_2554 + _GEN_2337; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2338 = {{3'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2556 = _T_2555 + _GEN_2338; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2339 = {{4'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2557 = _T_2556 + _GEN_2339; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2340 = {{5'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2558 = _T_2557 + _GEN_2340; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2341 = {{6'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2559 = _T_2558 + _GEN_2341; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2342 = {{7'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2560 = _T_2559 + _GEN_2342; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2343 = {{8'd0}, regs_10_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2562 = _T_2560 - _GEN_2343; // @[Conwaylife.scala 29:42]
  wire  _T_2563 = _T_2562 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2564 = _T_2562 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2565 = _T_2562 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2567 = regs_9_4 + regs_9_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2344 = {{1'd0}, regs_9_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2568 = _T_2567 + _GEN_2344; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2345 = {{2'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2569 = _T_2568 + _GEN_2345; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2346 = {{3'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2570 = _T_2569 + _GEN_2346; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2347 = {{4'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2571 = _T_2570 + _GEN_2347; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2348 = {{5'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2572 = _T_2571 + _GEN_2348; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2349 = {{6'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2573 = _T_2572 + _GEN_2349; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2350 = {{7'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2574 = _T_2573 + _GEN_2350; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2351 = {{8'd0}, regs_10_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2576 = _T_2574 - _GEN_2351; // @[Conwaylife.scala 29:42]
  wire  _T_2577 = _T_2576 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2578 = _T_2576 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2579 = _T_2576 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2581 = regs_9_5 + regs_9_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2352 = {{1'd0}, regs_9_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2582 = _T_2581 + _GEN_2352; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2353 = {{2'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2583 = _T_2582 + _GEN_2353; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2354 = {{3'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2584 = _T_2583 + _GEN_2354; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2355 = {{4'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2585 = _T_2584 + _GEN_2355; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2356 = {{5'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2586 = _T_2585 + _GEN_2356; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2357 = {{6'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2587 = _T_2586 + _GEN_2357; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2358 = {{7'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2588 = _T_2587 + _GEN_2358; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2359 = {{8'd0}, regs_10_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2590 = _T_2588 - _GEN_2359; // @[Conwaylife.scala 29:42]
  wire  _T_2591 = _T_2590 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2592 = _T_2590 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2593 = _T_2590 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2595 = regs_9_6 + regs_9_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2360 = {{1'd0}, regs_9_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2596 = _T_2595 + _GEN_2360; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2361 = {{2'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2597 = _T_2596 + _GEN_2361; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2362 = {{3'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2598 = _T_2597 + _GEN_2362; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2363 = {{4'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2599 = _T_2598 + _GEN_2363; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2364 = {{5'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2600 = _T_2599 + _GEN_2364; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2365 = {{6'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2601 = _T_2600 + _GEN_2365; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2366 = {{7'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2602 = _T_2601 + _GEN_2366; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2367 = {{8'd0}, regs_10_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2604 = _T_2602 - _GEN_2367; // @[Conwaylife.scala 29:42]
  wire  _T_2605 = _T_2604 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2606 = _T_2604 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2607 = _T_2604 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2609 = regs_9_7 + regs_9_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2368 = {{1'd0}, regs_9_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2610 = _T_2609 + _GEN_2368; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2369 = {{2'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2611 = _T_2610 + _GEN_2369; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2370 = {{3'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2612 = _T_2611 + _GEN_2370; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2371 = {{4'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2613 = _T_2612 + _GEN_2371; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2372 = {{5'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2614 = _T_2613 + _GEN_2372; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2373 = {{6'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2615 = _T_2614 + _GEN_2373; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2374 = {{7'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2616 = _T_2615 + _GEN_2374; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2375 = {{8'd0}, regs_10_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2618 = _T_2616 - _GEN_2375; // @[Conwaylife.scala 29:42]
  wire  _T_2619 = _T_2618 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2620 = _T_2618 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2621 = _T_2618 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2623 = regs_9_8 + regs_9_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2376 = {{1'd0}, regs_9_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2624 = _T_2623 + _GEN_2376; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2377 = {{2'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2625 = _T_2624 + _GEN_2377; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2378 = {{3'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2626 = _T_2625 + _GEN_2378; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2379 = {{4'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2627 = _T_2626 + _GEN_2379; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2380 = {{5'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2628 = _T_2627 + _GEN_2380; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2381 = {{6'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2629 = _T_2628 + _GEN_2381; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2382 = {{7'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2630 = _T_2629 + _GEN_2382; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2383 = {{8'd0}, regs_10_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2632 = _T_2630 - _GEN_2383; // @[Conwaylife.scala 29:42]
  wire  _T_2633 = _T_2632 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2634 = _T_2632 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2635 = _T_2632 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2637 = regs_9_9 + regs_9_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2384 = {{1'd0}, regs_9_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2638 = _T_2637 + _GEN_2384; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2385 = {{2'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2639 = _T_2638 + _GEN_2385; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2386 = {{3'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2640 = _T_2639 + _GEN_2386; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2387 = {{4'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2641 = _T_2640 + _GEN_2387; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2388 = {{5'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2642 = _T_2641 + _GEN_2388; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2389 = {{6'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2643 = _T_2642 + _GEN_2389; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2390 = {{7'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2644 = _T_2643 + _GEN_2390; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2391 = {{8'd0}, regs_10_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2646 = _T_2644 - _GEN_2391; // @[Conwaylife.scala 29:42]
  wire  _T_2647 = _T_2646 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2648 = _T_2646 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2649 = _T_2646 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2651 = regs_9_10 + regs_9_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2392 = {{1'd0}, regs_9_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2652 = _T_2651 + _GEN_2392; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2393 = {{2'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2653 = _T_2652 + _GEN_2393; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2394 = {{3'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2654 = _T_2653 + _GEN_2394; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2395 = {{4'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2655 = _T_2654 + _GEN_2395; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2396 = {{5'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2656 = _T_2655 + _GEN_2396; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2397 = {{6'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2657 = _T_2656 + _GEN_2397; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2398 = {{7'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2658 = _T_2657 + _GEN_2398; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2399 = {{8'd0}, regs_10_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2660 = _T_2658 - _GEN_2399; // @[Conwaylife.scala 29:42]
  wire  _T_2661 = _T_2660 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2662 = _T_2660 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2663 = _T_2660 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2665 = regs_9_11 + regs_9_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2400 = {{1'd0}, regs_9_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2666 = _T_2665 + _GEN_2400; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2401 = {{2'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2667 = _T_2666 + _GEN_2401; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2402 = {{3'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2668 = _T_2667 + _GEN_2402; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2403 = {{4'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2669 = _T_2668 + _GEN_2403; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2404 = {{5'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2670 = _T_2669 + _GEN_2404; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2405 = {{6'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2671 = _T_2670 + _GEN_2405; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2406 = {{7'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2672 = _T_2671 + _GEN_2406; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2407 = {{8'd0}, regs_10_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2674 = _T_2672 - _GEN_2407; // @[Conwaylife.scala 29:42]
  wire  _T_2675 = _T_2674 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2676 = _T_2674 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2677 = _T_2674 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2679 = regs_9_12 + regs_9_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2408 = {{1'd0}, regs_9_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2680 = _T_2679 + _GEN_2408; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2409 = {{2'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2681 = _T_2680 + _GEN_2409; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2410 = {{3'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2682 = _T_2681 + _GEN_2410; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2411 = {{4'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2683 = _T_2682 + _GEN_2411; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2412 = {{5'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2684 = _T_2683 + _GEN_2412; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2413 = {{6'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2685 = _T_2684 + _GEN_2413; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2414 = {{7'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2686 = _T_2685 + _GEN_2414; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2415 = {{8'd0}, regs_10_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2688 = _T_2686 - _GEN_2415; // @[Conwaylife.scala 29:42]
  wire  _T_2689 = _T_2688 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2690 = _T_2688 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2691 = _T_2688 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2693 = regs_9_13 + regs_9_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2416 = {{1'd0}, regs_9_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2694 = _T_2693 + _GEN_2416; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2417 = {{2'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2695 = _T_2694 + _GEN_2417; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2418 = {{3'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2696 = _T_2695 + _GEN_2418; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2419 = {{4'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2697 = _T_2696 + _GEN_2419; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2420 = {{5'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2698 = _T_2697 + _GEN_2420; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2421 = {{6'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2699 = _T_2698 + _GEN_2421; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2422 = {{7'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2700 = _T_2699 + _GEN_2422; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2423 = {{8'd0}, regs_10_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2702 = _T_2700 - _GEN_2423; // @[Conwaylife.scala 29:42]
  wire  _T_2703 = _T_2702 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2704 = _T_2702 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2705 = _T_2702 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2707 = regs_9_14 + regs_9_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2424 = {{1'd0}, regs_9_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2708 = _T_2707 + _GEN_2424; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2425 = {{2'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2709 = _T_2708 + _GEN_2425; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2426 = {{3'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2710 = _T_2709 + _GEN_2426; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2427 = {{4'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2711 = _T_2710 + _GEN_2427; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2428 = {{5'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2712 = _T_2711 + _GEN_2428; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2429 = {{6'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2713 = _T_2712 + _GEN_2429; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2430 = {{7'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2714 = _T_2713 + _GEN_2430; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2431 = {{8'd0}, regs_10_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2716 = _T_2714 - _GEN_2431; // @[Conwaylife.scala 29:42]
  wire  _T_2717 = _T_2716 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2718 = _T_2716 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2719 = _T_2716 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2721 = regs_10_15 + regs_10_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2432 = {{1'd0}, regs_10_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2722 = _T_2721 + _GEN_2432; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2433 = {{2'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2723 = _T_2722 + _GEN_2433; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2434 = {{3'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2724 = _T_2723 + _GEN_2434; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2435 = {{4'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2725 = _T_2724 + _GEN_2435; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2436 = {{5'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2726 = _T_2725 + _GEN_2436; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2437 = {{6'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2727 = _T_2726 + _GEN_2437; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2438 = {{7'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2728 = _T_2727 + _GEN_2438; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2439 = {{8'd0}, regs_11_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2730 = _T_2728 - _GEN_2439; // @[Conwaylife.scala 29:42]
  wire  _T_2731 = _T_2730 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2732 = _T_2730 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2733 = _T_2730 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2735 = regs_10_0 + regs_10_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2440 = {{1'd0}, regs_10_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2736 = _T_2735 + _GEN_2440; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2441 = {{2'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2737 = _T_2736 + _GEN_2441; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2442 = {{3'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2738 = _T_2737 + _GEN_2442; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2443 = {{4'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2739 = _T_2738 + _GEN_2443; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2444 = {{5'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2740 = _T_2739 + _GEN_2444; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2445 = {{6'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2741 = _T_2740 + _GEN_2445; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2446 = {{7'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2742 = _T_2741 + _GEN_2446; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2447 = {{8'd0}, regs_11_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2744 = _T_2742 - _GEN_2447; // @[Conwaylife.scala 29:42]
  wire  _T_2745 = _T_2744 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2746 = _T_2744 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2747 = _T_2744 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2749 = regs_10_1 + regs_10_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2448 = {{1'd0}, regs_10_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2750 = _T_2749 + _GEN_2448; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2449 = {{2'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2751 = _T_2750 + _GEN_2449; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2450 = {{3'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2752 = _T_2751 + _GEN_2450; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2451 = {{4'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2753 = _T_2752 + _GEN_2451; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2452 = {{5'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2754 = _T_2753 + _GEN_2452; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2453 = {{6'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2755 = _T_2754 + _GEN_2453; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2454 = {{7'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2756 = _T_2755 + _GEN_2454; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2455 = {{8'd0}, regs_11_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2758 = _T_2756 - _GEN_2455; // @[Conwaylife.scala 29:42]
  wire  _T_2759 = _T_2758 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2760 = _T_2758 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2761 = _T_2758 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2763 = regs_10_2 + regs_10_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2456 = {{1'd0}, regs_10_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2764 = _T_2763 + _GEN_2456; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2457 = {{2'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2765 = _T_2764 + _GEN_2457; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2458 = {{3'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2766 = _T_2765 + _GEN_2458; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2459 = {{4'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2767 = _T_2766 + _GEN_2459; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2460 = {{5'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2768 = _T_2767 + _GEN_2460; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2461 = {{6'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2769 = _T_2768 + _GEN_2461; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2462 = {{7'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2770 = _T_2769 + _GEN_2462; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2463 = {{8'd0}, regs_11_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2772 = _T_2770 - _GEN_2463; // @[Conwaylife.scala 29:42]
  wire  _T_2773 = _T_2772 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2774 = _T_2772 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2775 = _T_2772 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2777 = regs_10_3 + regs_10_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2464 = {{1'd0}, regs_10_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2778 = _T_2777 + _GEN_2464; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2465 = {{2'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2779 = _T_2778 + _GEN_2465; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2466 = {{3'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2780 = _T_2779 + _GEN_2466; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2467 = {{4'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2781 = _T_2780 + _GEN_2467; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2468 = {{5'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2782 = _T_2781 + _GEN_2468; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2469 = {{6'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2783 = _T_2782 + _GEN_2469; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2470 = {{7'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2784 = _T_2783 + _GEN_2470; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2471 = {{8'd0}, regs_11_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2786 = _T_2784 - _GEN_2471; // @[Conwaylife.scala 29:42]
  wire  _T_2787 = _T_2786 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2788 = _T_2786 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2789 = _T_2786 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2791 = regs_10_4 + regs_10_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2472 = {{1'd0}, regs_10_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2792 = _T_2791 + _GEN_2472; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2473 = {{2'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2793 = _T_2792 + _GEN_2473; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2474 = {{3'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2794 = _T_2793 + _GEN_2474; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2475 = {{4'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2795 = _T_2794 + _GEN_2475; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2476 = {{5'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2796 = _T_2795 + _GEN_2476; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2477 = {{6'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2797 = _T_2796 + _GEN_2477; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2478 = {{7'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2798 = _T_2797 + _GEN_2478; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2479 = {{8'd0}, regs_11_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2800 = _T_2798 - _GEN_2479; // @[Conwaylife.scala 29:42]
  wire  _T_2801 = _T_2800 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2802 = _T_2800 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2803 = _T_2800 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2805 = regs_10_5 + regs_10_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2480 = {{1'd0}, regs_10_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2806 = _T_2805 + _GEN_2480; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2481 = {{2'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2807 = _T_2806 + _GEN_2481; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2482 = {{3'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2808 = _T_2807 + _GEN_2482; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2483 = {{4'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2809 = _T_2808 + _GEN_2483; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2484 = {{5'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2810 = _T_2809 + _GEN_2484; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2485 = {{6'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2811 = _T_2810 + _GEN_2485; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2486 = {{7'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2812 = _T_2811 + _GEN_2486; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2487 = {{8'd0}, regs_11_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2814 = _T_2812 - _GEN_2487; // @[Conwaylife.scala 29:42]
  wire  _T_2815 = _T_2814 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2816 = _T_2814 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2817 = _T_2814 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2819 = regs_10_6 + regs_10_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2488 = {{1'd0}, regs_10_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2820 = _T_2819 + _GEN_2488; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2489 = {{2'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2821 = _T_2820 + _GEN_2489; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2490 = {{3'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2822 = _T_2821 + _GEN_2490; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2491 = {{4'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2823 = _T_2822 + _GEN_2491; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2492 = {{5'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2824 = _T_2823 + _GEN_2492; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2493 = {{6'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2825 = _T_2824 + _GEN_2493; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2494 = {{7'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2826 = _T_2825 + _GEN_2494; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2495 = {{8'd0}, regs_11_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2828 = _T_2826 - _GEN_2495; // @[Conwaylife.scala 29:42]
  wire  _T_2829 = _T_2828 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2830 = _T_2828 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2831 = _T_2828 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2833 = regs_10_7 + regs_10_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2496 = {{1'd0}, regs_10_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2834 = _T_2833 + _GEN_2496; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2497 = {{2'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2835 = _T_2834 + _GEN_2497; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2498 = {{3'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2836 = _T_2835 + _GEN_2498; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2499 = {{4'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2837 = _T_2836 + _GEN_2499; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2500 = {{5'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2838 = _T_2837 + _GEN_2500; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2501 = {{6'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2839 = _T_2838 + _GEN_2501; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2502 = {{7'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2840 = _T_2839 + _GEN_2502; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2503 = {{8'd0}, regs_11_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2842 = _T_2840 - _GEN_2503; // @[Conwaylife.scala 29:42]
  wire  _T_2843 = _T_2842 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2844 = _T_2842 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2845 = _T_2842 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2847 = regs_10_8 + regs_10_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2504 = {{1'd0}, regs_10_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2848 = _T_2847 + _GEN_2504; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2505 = {{2'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2849 = _T_2848 + _GEN_2505; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2506 = {{3'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2850 = _T_2849 + _GEN_2506; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2507 = {{4'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2851 = _T_2850 + _GEN_2507; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2508 = {{5'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2852 = _T_2851 + _GEN_2508; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2509 = {{6'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2853 = _T_2852 + _GEN_2509; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2510 = {{7'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2854 = _T_2853 + _GEN_2510; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2511 = {{8'd0}, regs_11_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2856 = _T_2854 - _GEN_2511; // @[Conwaylife.scala 29:42]
  wire  _T_2857 = _T_2856 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2858 = _T_2856 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2859 = _T_2856 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2861 = regs_10_9 + regs_10_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2512 = {{1'd0}, regs_10_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2862 = _T_2861 + _GEN_2512; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2513 = {{2'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2863 = _T_2862 + _GEN_2513; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2514 = {{3'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2864 = _T_2863 + _GEN_2514; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2515 = {{4'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2865 = _T_2864 + _GEN_2515; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2516 = {{5'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2866 = _T_2865 + _GEN_2516; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2517 = {{6'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2867 = _T_2866 + _GEN_2517; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2518 = {{7'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2868 = _T_2867 + _GEN_2518; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2519 = {{8'd0}, regs_11_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2870 = _T_2868 - _GEN_2519; // @[Conwaylife.scala 29:42]
  wire  _T_2871 = _T_2870 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2872 = _T_2870 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2873 = _T_2870 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2875 = regs_10_10 + regs_10_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2520 = {{1'd0}, regs_10_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2876 = _T_2875 + _GEN_2520; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2521 = {{2'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2877 = _T_2876 + _GEN_2521; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2522 = {{3'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2878 = _T_2877 + _GEN_2522; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2523 = {{4'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2879 = _T_2878 + _GEN_2523; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2524 = {{5'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2880 = _T_2879 + _GEN_2524; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2525 = {{6'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2881 = _T_2880 + _GEN_2525; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2526 = {{7'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2882 = _T_2881 + _GEN_2526; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2527 = {{8'd0}, regs_11_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2884 = _T_2882 - _GEN_2527; // @[Conwaylife.scala 29:42]
  wire  _T_2885 = _T_2884 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2886 = _T_2884 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2887 = _T_2884 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2889 = regs_10_11 + regs_10_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2528 = {{1'd0}, regs_10_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2890 = _T_2889 + _GEN_2528; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2529 = {{2'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2891 = _T_2890 + _GEN_2529; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2530 = {{3'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2892 = _T_2891 + _GEN_2530; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2531 = {{4'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2893 = _T_2892 + _GEN_2531; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2532 = {{5'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2894 = _T_2893 + _GEN_2532; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2533 = {{6'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2895 = _T_2894 + _GEN_2533; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2534 = {{7'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2896 = _T_2895 + _GEN_2534; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2535 = {{8'd0}, regs_11_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2898 = _T_2896 - _GEN_2535; // @[Conwaylife.scala 29:42]
  wire  _T_2899 = _T_2898 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2900 = _T_2898 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2901 = _T_2898 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2903 = regs_10_12 + regs_10_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2536 = {{1'd0}, regs_10_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2904 = _T_2903 + _GEN_2536; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2537 = {{2'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2905 = _T_2904 + _GEN_2537; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2538 = {{3'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2906 = _T_2905 + _GEN_2538; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2539 = {{4'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2907 = _T_2906 + _GEN_2539; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2540 = {{5'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2908 = _T_2907 + _GEN_2540; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2541 = {{6'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2909 = _T_2908 + _GEN_2541; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2542 = {{7'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2910 = _T_2909 + _GEN_2542; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2543 = {{8'd0}, regs_11_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2912 = _T_2910 - _GEN_2543; // @[Conwaylife.scala 29:42]
  wire  _T_2913 = _T_2912 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2914 = _T_2912 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2915 = _T_2912 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2917 = regs_10_13 + regs_10_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2544 = {{1'd0}, regs_10_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2918 = _T_2917 + _GEN_2544; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2545 = {{2'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2919 = _T_2918 + _GEN_2545; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2546 = {{3'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2920 = _T_2919 + _GEN_2546; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2547 = {{4'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2921 = _T_2920 + _GEN_2547; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2548 = {{5'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2922 = _T_2921 + _GEN_2548; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2549 = {{6'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2923 = _T_2922 + _GEN_2549; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2550 = {{7'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2924 = _T_2923 + _GEN_2550; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2551 = {{8'd0}, regs_11_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2926 = _T_2924 - _GEN_2551; // @[Conwaylife.scala 29:42]
  wire  _T_2927 = _T_2926 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2928 = _T_2926 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2929 = _T_2926 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2931 = regs_10_14 + regs_10_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2552 = {{1'd0}, regs_10_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2932 = _T_2931 + _GEN_2552; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2553 = {{2'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2933 = _T_2932 + _GEN_2553; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2554 = {{3'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2934 = _T_2933 + _GEN_2554; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2555 = {{4'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2935 = _T_2934 + _GEN_2555; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2556 = {{5'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2936 = _T_2935 + _GEN_2556; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2557 = {{6'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2937 = _T_2936 + _GEN_2557; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2558 = {{7'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2938 = _T_2937 + _GEN_2558; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2559 = {{8'd0}, regs_11_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2940 = _T_2938 - _GEN_2559; // @[Conwaylife.scala 29:42]
  wire  _T_2941 = _T_2940 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2942 = _T_2940 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2943 = _T_2940 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2945 = regs_11_15 + regs_11_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2560 = {{1'd0}, regs_11_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2946 = _T_2945 + _GEN_2560; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2561 = {{2'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2947 = _T_2946 + _GEN_2561; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2562 = {{3'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2948 = _T_2947 + _GEN_2562; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2563 = {{4'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2949 = _T_2948 + _GEN_2563; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2564 = {{5'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2950 = _T_2949 + _GEN_2564; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2565 = {{6'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2951 = _T_2950 + _GEN_2565; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2566 = {{7'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2952 = _T_2951 + _GEN_2566; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2567 = {{8'd0}, regs_12_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2954 = _T_2952 - _GEN_2567; // @[Conwaylife.scala 29:42]
  wire  _T_2955 = _T_2954 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2956 = _T_2954 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2957 = _T_2954 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2959 = regs_11_0 + regs_11_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2568 = {{1'd0}, regs_11_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2960 = _T_2959 + _GEN_2568; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2569 = {{2'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2961 = _T_2960 + _GEN_2569; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2570 = {{3'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2962 = _T_2961 + _GEN_2570; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2571 = {{4'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2963 = _T_2962 + _GEN_2571; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2572 = {{5'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2964 = _T_2963 + _GEN_2572; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2573 = {{6'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2965 = _T_2964 + _GEN_2573; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2574 = {{7'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2966 = _T_2965 + _GEN_2574; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2575 = {{8'd0}, regs_12_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2968 = _T_2966 - _GEN_2575; // @[Conwaylife.scala 29:42]
  wire  _T_2969 = _T_2968 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2970 = _T_2968 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2971 = _T_2968 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2973 = regs_11_1 + regs_11_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2576 = {{1'd0}, regs_11_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2974 = _T_2973 + _GEN_2576; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2577 = {{2'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2975 = _T_2974 + _GEN_2577; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2578 = {{3'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2976 = _T_2975 + _GEN_2578; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2579 = {{4'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2977 = _T_2976 + _GEN_2579; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2580 = {{5'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2978 = _T_2977 + _GEN_2580; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2581 = {{6'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2979 = _T_2978 + _GEN_2581; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2582 = {{7'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2980 = _T_2979 + _GEN_2582; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2583 = {{8'd0}, regs_12_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2982 = _T_2980 - _GEN_2583; // @[Conwaylife.scala 29:42]
  wire  _T_2983 = _T_2982 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2984 = _T_2982 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2985 = _T_2982 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_2987 = regs_11_2 + regs_11_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2584 = {{1'd0}, regs_11_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_2988 = _T_2987 + _GEN_2584; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2585 = {{2'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_2989 = _T_2988 + _GEN_2585; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2586 = {{3'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_2990 = _T_2989 + _GEN_2586; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2587 = {{4'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_2991 = _T_2990 + _GEN_2587; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2588 = {{5'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_2992 = _T_2991 + _GEN_2588; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2589 = {{6'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_2993 = _T_2992 + _GEN_2589; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2590 = {{7'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_2994 = _T_2993 + _GEN_2590; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2591 = {{8'd0}, regs_12_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_2996 = _T_2994 - _GEN_2591; // @[Conwaylife.scala 29:42]
  wire  _T_2997 = _T_2996 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_2998 = _T_2996 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_2999 = _T_2996 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3001 = regs_11_3 + regs_11_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2592 = {{1'd0}, regs_11_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3002 = _T_3001 + _GEN_2592; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2593 = {{2'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3003 = _T_3002 + _GEN_2593; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2594 = {{3'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3004 = _T_3003 + _GEN_2594; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2595 = {{4'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3005 = _T_3004 + _GEN_2595; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2596 = {{5'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3006 = _T_3005 + _GEN_2596; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2597 = {{6'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3007 = _T_3006 + _GEN_2597; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2598 = {{7'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3008 = _T_3007 + _GEN_2598; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2599 = {{8'd0}, regs_12_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3010 = _T_3008 - _GEN_2599; // @[Conwaylife.scala 29:42]
  wire  _T_3011 = _T_3010 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3012 = _T_3010 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3013 = _T_3010 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3015 = regs_11_4 + regs_11_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2600 = {{1'd0}, regs_11_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3016 = _T_3015 + _GEN_2600; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2601 = {{2'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3017 = _T_3016 + _GEN_2601; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2602 = {{3'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3018 = _T_3017 + _GEN_2602; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2603 = {{4'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3019 = _T_3018 + _GEN_2603; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2604 = {{5'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3020 = _T_3019 + _GEN_2604; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2605 = {{6'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3021 = _T_3020 + _GEN_2605; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2606 = {{7'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3022 = _T_3021 + _GEN_2606; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2607 = {{8'd0}, regs_12_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3024 = _T_3022 - _GEN_2607; // @[Conwaylife.scala 29:42]
  wire  _T_3025 = _T_3024 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3026 = _T_3024 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3027 = _T_3024 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3029 = regs_11_5 + regs_11_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2608 = {{1'd0}, regs_11_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3030 = _T_3029 + _GEN_2608; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2609 = {{2'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3031 = _T_3030 + _GEN_2609; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2610 = {{3'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3032 = _T_3031 + _GEN_2610; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2611 = {{4'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3033 = _T_3032 + _GEN_2611; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2612 = {{5'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3034 = _T_3033 + _GEN_2612; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2613 = {{6'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3035 = _T_3034 + _GEN_2613; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2614 = {{7'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3036 = _T_3035 + _GEN_2614; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2615 = {{8'd0}, regs_12_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3038 = _T_3036 - _GEN_2615; // @[Conwaylife.scala 29:42]
  wire  _T_3039 = _T_3038 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3040 = _T_3038 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3041 = _T_3038 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3043 = regs_11_6 + regs_11_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2616 = {{1'd0}, regs_11_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3044 = _T_3043 + _GEN_2616; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2617 = {{2'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3045 = _T_3044 + _GEN_2617; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2618 = {{3'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3046 = _T_3045 + _GEN_2618; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2619 = {{4'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3047 = _T_3046 + _GEN_2619; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2620 = {{5'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3048 = _T_3047 + _GEN_2620; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2621 = {{6'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3049 = _T_3048 + _GEN_2621; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2622 = {{7'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3050 = _T_3049 + _GEN_2622; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2623 = {{8'd0}, regs_12_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3052 = _T_3050 - _GEN_2623; // @[Conwaylife.scala 29:42]
  wire  _T_3053 = _T_3052 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3054 = _T_3052 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3055 = _T_3052 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3057 = regs_11_7 + regs_11_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2624 = {{1'd0}, regs_11_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3058 = _T_3057 + _GEN_2624; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2625 = {{2'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3059 = _T_3058 + _GEN_2625; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2626 = {{3'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3060 = _T_3059 + _GEN_2626; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2627 = {{4'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3061 = _T_3060 + _GEN_2627; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2628 = {{5'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3062 = _T_3061 + _GEN_2628; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2629 = {{6'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3063 = _T_3062 + _GEN_2629; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2630 = {{7'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3064 = _T_3063 + _GEN_2630; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2631 = {{8'd0}, regs_12_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3066 = _T_3064 - _GEN_2631; // @[Conwaylife.scala 29:42]
  wire  _T_3067 = _T_3066 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3068 = _T_3066 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3069 = _T_3066 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3071 = regs_11_8 + regs_11_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2632 = {{1'd0}, regs_11_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3072 = _T_3071 + _GEN_2632; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2633 = {{2'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3073 = _T_3072 + _GEN_2633; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2634 = {{3'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3074 = _T_3073 + _GEN_2634; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2635 = {{4'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3075 = _T_3074 + _GEN_2635; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2636 = {{5'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3076 = _T_3075 + _GEN_2636; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2637 = {{6'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3077 = _T_3076 + _GEN_2637; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2638 = {{7'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3078 = _T_3077 + _GEN_2638; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2639 = {{8'd0}, regs_12_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3080 = _T_3078 - _GEN_2639; // @[Conwaylife.scala 29:42]
  wire  _T_3081 = _T_3080 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3082 = _T_3080 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3083 = _T_3080 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3085 = regs_11_9 + regs_11_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2640 = {{1'd0}, regs_11_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3086 = _T_3085 + _GEN_2640; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2641 = {{2'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3087 = _T_3086 + _GEN_2641; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2642 = {{3'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3088 = _T_3087 + _GEN_2642; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2643 = {{4'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3089 = _T_3088 + _GEN_2643; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2644 = {{5'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3090 = _T_3089 + _GEN_2644; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2645 = {{6'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3091 = _T_3090 + _GEN_2645; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2646 = {{7'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3092 = _T_3091 + _GEN_2646; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2647 = {{8'd0}, regs_12_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3094 = _T_3092 - _GEN_2647; // @[Conwaylife.scala 29:42]
  wire  _T_3095 = _T_3094 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3096 = _T_3094 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3097 = _T_3094 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3099 = regs_11_10 + regs_11_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2648 = {{1'd0}, regs_11_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3100 = _T_3099 + _GEN_2648; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2649 = {{2'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3101 = _T_3100 + _GEN_2649; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2650 = {{3'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3102 = _T_3101 + _GEN_2650; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2651 = {{4'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3103 = _T_3102 + _GEN_2651; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2652 = {{5'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3104 = _T_3103 + _GEN_2652; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2653 = {{6'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3105 = _T_3104 + _GEN_2653; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2654 = {{7'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3106 = _T_3105 + _GEN_2654; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2655 = {{8'd0}, regs_12_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3108 = _T_3106 - _GEN_2655; // @[Conwaylife.scala 29:42]
  wire  _T_3109 = _T_3108 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3110 = _T_3108 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3111 = _T_3108 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3113 = regs_11_11 + regs_11_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2656 = {{1'd0}, regs_11_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3114 = _T_3113 + _GEN_2656; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2657 = {{2'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3115 = _T_3114 + _GEN_2657; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2658 = {{3'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3116 = _T_3115 + _GEN_2658; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2659 = {{4'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3117 = _T_3116 + _GEN_2659; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2660 = {{5'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3118 = _T_3117 + _GEN_2660; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2661 = {{6'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3119 = _T_3118 + _GEN_2661; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2662 = {{7'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3120 = _T_3119 + _GEN_2662; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2663 = {{8'd0}, regs_12_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3122 = _T_3120 - _GEN_2663; // @[Conwaylife.scala 29:42]
  wire  _T_3123 = _T_3122 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3124 = _T_3122 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3125 = _T_3122 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3127 = regs_11_12 + regs_11_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2664 = {{1'd0}, regs_11_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3128 = _T_3127 + _GEN_2664; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2665 = {{2'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3129 = _T_3128 + _GEN_2665; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2666 = {{3'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3130 = _T_3129 + _GEN_2666; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2667 = {{4'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3131 = _T_3130 + _GEN_2667; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2668 = {{5'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3132 = _T_3131 + _GEN_2668; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2669 = {{6'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3133 = _T_3132 + _GEN_2669; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2670 = {{7'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3134 = _T_3133 + _GEN_2670; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2671 = {{8'd0}, regs_12_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3136 = _T_3134 - _GEN_2671; // @[Conwaylife.scala 29:42]
  wire  _T_3137 = _T_3136 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3138 = _T_3136 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3139 = _T_3136 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3141 = regs_11_13 + regs_11_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2672 = {{1'd0}, regs_11_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3142 = _T_3141 + _GEN_2672; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2673 = {{2'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3143 = _T_3142 + _GEN_2673; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2674 = {{3'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3144 = _T_3143 + _GEN_2674; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2675 = {{4'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3145 = _T_3144 + _GEN_2675; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2676 = {{5'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3146 = _T_3145 + _GEN_2676; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2677 = {{6'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3147 = _T_3146 + _GEN_2677; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2678 = {{7'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3148 = _T_3147 + _GEN_2678; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2679 = {{8'd0}, regs_12_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3150 = _T_3148 - _GEN_2679; // @[Conwaylife.scala 29:42]
  wire  _T_3151 = _T_3150 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3152 = _T_3150 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3153 = _T_3150 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3155 = regs_11_14 + regs_11_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2680 = {{1'd0}, regs_11_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3156 = _T_3155 + _GEN_2680; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2681 = {{2'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3157 = _T_3156 + _GEN_2681; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2682 = {{3'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3158 = _T_3157 + _GEN_2682; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2683 = {{4'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3159 = _T_3158 + _GEN_2683; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2684 = {{5'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3160 = _T_3159 + _GEN_2684; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2685 = {{6'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3161 = _T_3160 + _GEN_2685; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2686 = {{7'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3162 = _T_3161 + _GEN_2686; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2687 = {{8'd0}, regs_12_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3164 = _T_3162 - _GEN_2687; // @[Conwaylife.scala 29:42]
  wire  _T_3165 = _T_3164 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3166 = _T_3164 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3167 = _T_3164 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3169 = regs_12_15 + regs_12_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2688 = {{1'd0}, regs_12_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3170 = _T_3169 + _GEN_2688; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2689 = {{2'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3171 = _T_3170 + _GEN_2689; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2690 = {{3'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3172 = _T_3171 + _GEN_2690; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2691 = {{4'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3173 = _T_3172 + _GEN_2691; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2692 = {{5'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3174 = _T_3173 + _GEN_2692; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2693 = {{6'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3175 = _T_3174 + _GEN_2693; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2694 = {{7'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3176 = _T_3175 + _GEN_2694; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2695 = {{8'd0}, regs_13_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3178 = _T_3176 - _GEN_2695; // @[Conwaylife.scala 29:42]
  wire  _T_3179 = _T_3178 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3180 = _T_3178 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3181 = _T_3178 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3183 = regs_12_0 + regs_12_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2696 = {{1'd0}, regs_12_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3184 = _T_3183 + _GEN_2696; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2697 = {{2'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3185 = _T_3184 + _GEN_2697; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2698 = {{3'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3186 = _T_3185 + _GEN_2698; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2699 = {{4'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3187 = _T_3186 + _GEN_2699; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2700 = {{5'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3188 = _T_3187 + _GEN_2700; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2701 = {{6'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3189 = _T_3188 + _GEN_2701; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2702 = {{7'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3190 = _T_3189 + _GEN_2702; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2703 = {{8'd0}, regs_13_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3192 = _T_3190 - _GEN_2703; // @[Conwaylife.scala 29:42]
  wire  _T_3193 = _T_3192 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3194 = _T_3192 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3195 = _T_3192 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3197 = regs_12_1 + regs_12_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2704 = {{1'd0}, regs_12_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3198 = _T_3197 + _GEN_2704; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2705 = {{2'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3199 = _T_3198 + _GEN_2705; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2706 = {{3'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3200 = _T_3199 + _GEN_2706; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2707 = {{4'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3201 = _T_3200 + _GEN_2707; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2708 = {{5'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3202 = _T_3201 + _GEN_2708; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2709 = {{6'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3203 = _T_3202 + _GEN_2709; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2710 = {{7'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3204 = _T_3203 + _GEN_2710; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2711 = {{8'd0}, regs_13_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3206 = _T_3204 - _GEN_2711; // @[Conwaylife.scala 29:42]
  wire  _T_3207 = _T_3206 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3208 = _T_3206 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3209 = _T_3206 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3211 = regs_12_2 + regs_12_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2712 = {{1'd0}, regs_12_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3212 = _T_3211 + _GEN_2712; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2713 = {{2'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3213 = _T_3212 + _GEN_2713; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2714 = {{3'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3214 = _T_3213 + _GEN_2714; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2715 = {{4'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3215 = _T_3214 + _GEN_2715; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2716 = {{5'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3216 = _T_3215 + _GEN_2716; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2717 = {{6'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3217 = _T_3216 + _GEN_2717; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2718 = {{7'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3218 = _T_3217 + _GEN_2718; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2719 = {{8'd0}, regs_13_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3220 = _T_3218 - _GEN_2719; // @[Conwaylife.scala 29:42]
  wire  _T_3221 = _T_3220 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3222 = _T_3220 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3223 = _T_3220 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3225 = regs_12_3 + regs_12_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2720 = {{1'd0}, regs_12_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3226 = _T_3225 + _GEN_2720; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2721 = {{2'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3227 = _T_3226 + _GEN_2721; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2722 = {{3'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3228 = _T_3227 + _GEN_2722; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2723 = {{4'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3229 = _T_3228 + _GEN_2723; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2724 = {{5'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3230 = _T_3229 + _GEN_2724; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2725 = {{6'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3231 = _T_3230 + _GEN_2725; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2726 = {{7'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3232 = _T_3231 + _GEN_2726; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2727 = {{8'd0}, regs_13_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3234 = _T_3232 - _GEN_2727; // @[Conwaylife.scala 29:42]
  wire  _T_3235 = _T_3234 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3236 = _T_3234 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3237 = _T_3234 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3239 = regs_12_4 + regs_12_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2728 = {{1'd0}, regs_12_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3240 = _T_3239 + _GEN_2728; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2729 = {{2'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3241 = _T_3240 + _GEN_2729; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2730 = {{3'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3242 = _T_3241 + _GEN_2730; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2731 = {{4'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3243 = _T_3242 + _GEN_2731; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2732 = {{5'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3244 = _T_3243 + _GEN_2732; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2733 = {{6'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3245 = _T_3244 + _GEN_2733; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2734 = {{7'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3246 = _T_3245 + _GEN_2734; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2735 = {{8'd0}, regs_13_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3248 = _T_3246 - _GEN_2735; // @[Conwaylife.scala 29:42]
  wire  _T_3249 = _T_3248 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3250 = _T_3248 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3251 = _T_3248 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3253 = regs_12_5 + regs_12_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2736 = {{1'd0}, regs_12_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3254 = _T_3253 + _GEN_2736; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2737 = {{2'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3255 = _T_3254 + _GEN_2737; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2738 = {{3'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3256 = _T_3255 + _GEN_2738; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2739 = {{4'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3257 = _T_3256 + _GEN_2739; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2740 = {{5'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3258 = _T_3257 + _GEN_2740; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2741 = {{6'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3259 = _T_3258 + _GEN_2741; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2742 = {{7'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3260 = _T_3259 + _GEN_2742; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2743 = {{8'd0}, regs_13_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3262 = _T_3260 - _GEN_2743; // @[Conwaylife.scala 29:42]
  wire  _T_3263 = _T_3262 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3264 = _T_3262 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3265 = _T_3262 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3267 = regs_12_6 + regs_12_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2744 = {{1'd0}, regs_12_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3268 = _T_3267 + _GEN_2744; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2745 = {{2'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3269 = _T_3268 + _GEN_2745; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2746 = {{3'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3270 = _T_3269 + _GEN_2746; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2747 = {{4'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3271 = _T_3270 + _GEN_2747; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2748 = {{5'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3272 = _T_3271 + _GEN_2748; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2749 = {{6'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3273 = _T_3272 + _GEN_2749; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2750 = {{7'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3274 = _T_3273 + _GEN_2750; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2751 = {{8'd0}, regs_13_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3276 = _T_3274 - _GEN_2751; // @[Conwaylife.scala 29:42]
  wire  _T_3277 = _T_3276 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3278 = _T_3276 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3279 = _T_3276 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3281 = regs_12_7 + regs_12_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2752 = {{1'd0}, regs_12_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3282 = _T_3281 + _GEN_2752; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2753 = {{2'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3283 = _T_3282 + _GEN_2753; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2754 = {{3'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3284 = _T_3283 + _GEN_2754; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2755 = {{4'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3285 = _T_3284 + _GEN_2755; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2756 = {{5'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3286 = _T_3285 + _GEN_2756; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2757 = {{6'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3287 = _T_3286 + _GEN_2757; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2758 = {{7'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3288 = _T_3287 + _GEN_2758; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2759 = {{8'd0}, regs_13_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3290 = _T_3288 - _GEN_2759; // @[Conwaylife.scala 29:42]
  wire  _T_3291 = _T_3290 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3292 = _T_3290 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3293 = _T_3290 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3295 = regs_12_8 + regs_12_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2760 = {{1'd0}, regs_12_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3296 = _T_3295 + _GEN_2760; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2761 = {{2'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3297 = _T_3296 + _GEN_2761; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2762 = {{3'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3298 = _T_3297 + _GEN_2762; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2763 = {{4'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3299 = _T_3298 + _GEN_2763; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2764 = {{5'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3300 = _T_3299 + _GEN_2764; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2765 = {{6'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3301 = _T_3300 + _GEN_2765; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2766 = {{7'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3302 = _T_3301 + _GEN_2766; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2767 = {{8'd0}, regs_13_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3304 = _T_3302 - _GEN_2767; // @[Conwaylife.scala 29:42]
  wire  _T_3305 = _T_3304 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3306 = _T_3304 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3307 = _T_3304 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3309 = regs_12_9 + regs_12_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2768 = {{1'd0}, regs_12_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3310 = _T_3309 + _GEN_2768; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2769 = {{2'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3311 = _T_3310 + _GEN_2769; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2770 = {{3'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3312 = _T_3311 + _GEN_2770; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2771 = {{4'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3313 = _T_3312 + _GEN_2771; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2772 = {{5'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3314 = _T_3313 + _GEN_2772; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2773 = {{6'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3315 = _T_3314 + _GEN_2773; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2774 = {{7'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3316 = _T_3315 + _GEN_2774; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2775 = {{8'd0}, regs_13_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3318 = _T_3316 - _GEN_2775; // @[Conwaylife.scala 29:42]
  wire  _T_3319 = _T_3318 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3320 = _T_3318 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3321 = _T_3318 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3323 = regs_12_10 + regs_12_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2776 = {{1'd0}, regs_12_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3324 = _T_3323 + _GEN_2776; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2777 = {{2'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3325 = _T_3324 + _GEN_2777; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2778 = {{3'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3326 = _T_3325 + _GEN_2778; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2779 = {{4'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3327 = _T_3326 + _GEN_2779; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2780 = {{5'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3328 = _T_3327 + _GEN_2780; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2781 = {{6'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3329 = _T_3328 + _GEN_2781; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2782 = {{7'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3330 = _T_3329 + _GEN_2782; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2783 = {{8'd0}, regs_13_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3332 = _T_3330 - _GEN_2783; // @[Conwaylife.scala 29:42]
  wire  _T_3333 = _T_3332 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3334 = _T_3332 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3335 = _T_3332 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3337 = regs_12_11 + regs_12_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2784 = {{1'd0}, regs_12_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3338 = _T_3337 + _GEN_2784; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2785 = {{2'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3339 = _T_3338 + _GEN_2785; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2786 = {{3'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3340 = _T_3339 + _GEN_2786; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2787 = {{4'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3341 = _T_3340 + _GEN_2787; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2788 = {{5'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3342 = _T_3341 + _GEN_2788; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2789 = {{6'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3343 = _T_3342 + _GEN_2789; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2790 = {{7'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3344 = _T_3343 + _GEN_2790; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2791 = {{8'd0}, regs_13_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3346 = _T_3344 - _GEN_2791; // @[Conwaylife.scala 29:42]
  wire  _T_3347 = _T_3346 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3348 = _T_3346 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3349 = _T_3346 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3351 = regs_12_12 + regs_12_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2792 = {{1'd0}, regs_12_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3352 = _T_3351 + _GEN_2792; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2793 = {{2'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3353 = _T_3352 + _GEN_2793; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2794 = {{3'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3354 = _T_3353 + _GEN_2794; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2795 = {{4'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3355 = _T_3354 + _GEN_2795; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2796 = {{5'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3356 = _T_3355 + _GEN_2796; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2797 = {{6'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3357 = _T_3356 + _GEN_2797; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2798 = {{7'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3358 = _T_3357 + _GEN_2798; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2799 = {{8'd0}, regs_13_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3360 = _T_3358 - _GEN_2799; // @[Conwaylife.scala 29:42]
  wire  _T_3361 = _T_3360 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3362 = _T_3360 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3363 = _T_3360 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3365 = regs_12_13 + regs_12_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2800 = {{1'd0}, regs_12_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3366 = _T_3365 + _GEN_2800; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2801 = {{2'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3367 = _T_3366 + _GEN_2801; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2802 = {{3'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3368 = _T_3367 + _GEN_2802; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2803 = {{4'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3369 = _T_3368 + _GEN_2803; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2804 = {{5'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3370 = _T_3369 + _GEN_2804; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2805 = {{6'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3371 = _T_3370 + _GEN_2805; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2806 = {{7'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3372 = _T_3371 + _GEN_2806; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2807 = {{8'd0}, regs_13_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3374 = _T_3372 - _GEN_2807; // @[Conwaylife.scala 29:42]
  wire  _T_3375 = _T_3374 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3376 = _T_3374 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3377 = _T_3374 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3379 = regs_12_14 + regs_12_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2808 = {{1'd0}, regs_12_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3380 = _T_3379 + _GEN_2808; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2809 = {{2'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3381 = _T_3380 + _GEN_2809; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2810 = {{3'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3382 = _T_3381 + _GEN_2810; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2811 = {{4'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3383 = _T_3382 + _GEN_2811; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2812 = {{5'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3384 = _T_3383 + _GEN_2812; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2813 = {{6'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3385 = _T_3384 + _GEN_2813; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2814 = {{7'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3386 = _T_3385 + _GEN_2814; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2815 = {{8'd0}, regs_13_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3388 = _T_3386 - _GEN_2815; // @[Conwaylife.scala 29:42]
  wire  _T_3389 = _T_3388 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3390 = _T_3388 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3391 = _T_3388 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3393 = regs_13_15 + regs_13_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2816 = {{1'd0}, regs_13_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3394 = _T_3393 + _GEN_2816; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2817 = {{2'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3395 = _T_3394 + _GEN_2817; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2818 = {{3'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3396 = _T_3395 + _GEN_2818; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2819 = {{4'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3397 = _T_3396 + _GEN_2819; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2820 = {{5'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3398 = _T_3397 + _GEN_2820; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2821 = {{6'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3399 = _T_3398 + _GEN_2821; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2822 = {{7'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3400 = _T_3399 + _GEN_2822; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2823 = {{8'd0}, regs_14_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3402 = _T_3400 - _GEN_2823; // @[Conwaylife.scala 29:42]
  wire  _T_3403 = _T_3402 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3404 = _T_3402 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3405 = _T_3402 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3407 = regs_13_0 + regs_13_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2824 = {{1'd0}, regs_13_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3408 = _T_3407 + _GEN_2824; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2825 = {{2'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3409 = _T_3408 + _GEN_2825; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2826 = {{3'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3410 = _T_3409 + _GEN_2826; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2827 = {{4'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3411 = _T_3410 + _GEN_2827; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2828 = {{5'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3412 = _T_3411 + _GEN_2828; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2829 = {{6'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3413 = _T_3412 + _GEN_2829; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2830 = {{7'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3414 = _T_3413 + _GEN_2830; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2831 = {{8'd0}, regs_14_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3416 = _T_3414 - _GEN_2831; // @[Conwaylife.scala 29:42]
  wire  _T_3417 = _T_3416 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3418 = _T_3416 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3419 = _T_3416 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3421 = regs_13_1 + regs_13_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2832 = {{1'd0}, regs_13_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3422 = _T_3421 + _GEN_2832; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2833 = {{2'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3423 = _T_3422 + _GEN_2833; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2834 = {{3'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3424 = _T_3423 + _GEN_2834; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2835 = {{4'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3425 = _T_3424 + _GEN_2835; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2836 = {{5'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3426 = _T_3425 + _GEN_2836; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2837 = {{6'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3427 = _T_3426 + _GEN_2837; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2838 = {{7'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3428 = _T_3427 + _GEN_2838; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2839 = {{8'd0}, regs_14_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3430 = _T_3428 - _GEN_2839; // @[Conwaylife.scala 29:42]
  wire  _T_3431 = _T_3430 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3432 = _T_3430 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3433 = _T_3430 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3435 = regs_13_2 + regs_13_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2840 = {{1'd0}, regs_13_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3436 = _T_3435 + _GEN_2840; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2841 = {{2'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3437 = _T_3436 + _GEN_2841; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2842 = {{3'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3438 = _T_3437 + _GEN_2842; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2843 = {{4'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3439 = _T_3438 + _GEN_2843; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2844 = {{5'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3440 = _T_3439 + _GEN_2844; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2845 = {{6'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3441 = _T_3440 + _GEN_2845; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2846 = {{7'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3442 = _T_3441 + _GEN_2846; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2847 = {{8'd0}, regs_14_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3444 = _T_3442 - _GEN_2847; // @[Conwaylife.scala 29:42]
  wire  _T_3445 = _T_3444 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3446 = _T_3444 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3447 = _T_3444 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3449 = regs_13_3 + regs_13_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2848 = {{1'd0}, regs_13_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3450 = _T_3449 + _GEN_2848; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2849 = {{2'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3451 = _T_3450 + _GEN_2849; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2850 = {{3'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3452 = _T_3451 + _GEN_2850; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2851 = {{4'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3453 = _T_3452 + _GEN_2851; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2852 = {{5'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3454 = _T_3453 + _GEN_2852; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2853 = {{6'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3455 = _T_3454 + _GEN_2853; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2854 = {{7'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3456 = _T_3455 + _GEN_2854; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2855 = {{8'd0}, regs_14_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3458 = _T_3456 - _GEN_2855; // @[Conwaylife.scala 29:42]
  wire  _T_3459 = _T_3458 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3460 = _T_3458 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3461 = _T_3458 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3463 = regs_13_4 + regs_13_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2856 = {{1'd0}, regs_13_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3464 = _T_3463 + _GEN_2856; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2857 = {{2'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3465 = _T_3464 + _GEN_2857; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2858 = {{3'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3466 = _T_3465 + _GEN_2858; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2859 = {{4'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3467 = _T_3466 + _GEN_2859; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2860 = {{5'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3468 = _T_3467 + _GEN_2860; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2861 = {{6'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3469 = _T_3468 + _GEN_2861; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2862 = {{7'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3470 = _T_3469 + _GEN_2862; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2863 = {{8'd0}, regs_14_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3472 = _T_3470 - _GEN_2863; // @[Conwaylife.scala 29:42]
  wire  _T_3473 = _T_3472 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3474 = _T_3472 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3475 = _T_3472 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3477 = regs_13_5 + regs_13_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2864 = {{1'd0}, regs_13_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3478 = _T_3477 + _GEN_2864; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2865 = {{2'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3479 = _T_3478 + _GEN_2865; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2866 = {{3'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3480 = _T_3479 + _GEN_2866; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2867 = {{4'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3481 = _T_3480 + _GEN_2867; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2868 = {{5'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3482 = _T_3481 + _GEN_2868; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2869 = {{6'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3483 = _T_3482 + _GEN_2869; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2870 = {{7'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3484 = _T_3483 + _GEN_2870; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2871 = {{8'd0}, regs_14_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3486 = _T_3484 - _GEN_2871; // @[Conwaylife.scala 29:42]
  wire  _T_3487 = _T_3486 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3488 = _T_3486 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3489 = _T_3486 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3491 = regs_13_6 + regs_13_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2872 = {{1'd0}, regs_13_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3492 = _T_3491 + _GEN_2872; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2873 = {{2'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3493 = _T_3492 + _GEN_2873; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2874 = {{3'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3494 = _T_3493 + _GEN_2874; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2875 = {{4'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3495 = _T_3494 + _GEN_2875; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2876 = {{5'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3496 = _T_3495 + _GEN_2876; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2877 = {{6'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3497 = _T_3496 + _GEN_2877; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2878 = {{7'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3498 = _T_3497 + _GEN_2878; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2879 = {{8'd0}, regs_14_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3500 = _T_3498 - _GEN_2879; // @[Conwaylife.scala 29:42]
  wire  _T_3501 = _T_3500 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3502 = _T_3500 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3503 = _T_3500 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3505 = regs_13_7 + regs_13_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2880 = {{1'd0}, regs_13_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3506 = _T_3505 + _GEN_2880; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2881 = {{2'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3507 = _T_3506 + _GEN_2881; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2882 = {{3'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3508 = _T_3507 + _GEN_2882; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2883 = {{4'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3509 = _T_3508 + _GEN_2883; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2884 = {{5'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3510 = _T_3509 + _GEN_2884; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2885 = {{6'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3511 = _T_3510 + _GEN_2885; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2886 = {{7'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3512 = _T_3511 + _GEN_2886; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2887 = {{8'd0}, regs_14_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3514 = _T_3512 - _GEN_2887; // @[Conwaylife.scala 29:42]
  wire  _T_3515 = _T_3514 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3516 = _T_3514 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3517 = _T_3514 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3519 = regs_13_8 + regs_13_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2888 = {{1'd0}, regs_13_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3520 = _T_3519 + _GEN_2888; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2889 = {{2'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3521 = _T_3520 + _GEN_2889; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2890 = {{3'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3522 = _T_3521 + _GEN_2890; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2891 = {{4'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3523 = _T_3522 + _GEN_2891; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2892 = {{5'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3524 = _T_3523 + _GEN_2892; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2893 = {{6'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3525 = _T_3524 + _GEN_2893; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2894 = {{7'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3526 = _T_3525 + _GEN_2894; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2895 = {{8'd0}, regs_14_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3528 = _T_3526 - _GEN_2895; // @[Conwaylife.scala 29:42]
  wire  _T_3529 = _T_3528 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3530 = _T_3528 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3531 = _T_3528 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3533 = regs_13_9 + regs_13_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2896 = {{1'd0}, regs_13_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3534 = _T_3533 + _GEN_2896; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2897 = {{2'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3535 = _T_3534 + _GEN_2897; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2898 = {{3'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3536 = _T_3535 + _GEN_2898; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2899 = {{4'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3537 = _T_3536 + _GEN_2899; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2900 = {{5'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3538 = _T_3537 + _GEN_2900; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2901 = {{6'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3539 = _T_3538 + _GEN_2901; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2902 = {{7'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3540 = _T_3539 + _GEN_2902; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2903 = {{8'd0}, regs_14_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3542 = _T_3540 - _GEN_2903; // @[Conwaylife.scala 29:42]
  wire  _T_3543 = _T_3542 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3544 = _T_3542 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3545 = _T_3542 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3547 = regs_13_10 + regs_13_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2904 = {{1'd0}, regs_13_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3548 = _T_3547 + _GEN_2904; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2905 = {{2'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3549 = _T_3548 + _GEN_2905; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2906 = {{3'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3550 = _T_3549 + _GEN_2906; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2907 = {{4'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3551 = _T_3550 + _GEN_2907; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2908 = {{5'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3552 = _T_3551 + _GEN_2908; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2909 = {{6'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3553 = _T_3552 + _GEN_2909; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2910 = {{7'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3554 = _T_3553 + _GEN_2910; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2911 = {{8'd0}, regs_14_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3556 = _T_3554 - _GEN_2911; // @[Conwaylife.scala 29:42]
  wire  _T_3557 = _T_3556 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3558 = _T_3556 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3559 = _T_3556 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3561 = regs_13_11 + regs_13_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2912 = {{1'd0}, regs_13_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3562 = _T_3561 + _GEN_2912; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2913 = {{2'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3563 = _T_3562 + _GEN_2913; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2914 = {{3'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3564 = _T_3563 + _GEN_2914; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2915 = {{4'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3565 = _T_3564 + _GEN_2915; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2916 = {{5'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3566 = _T_3565 + _GEN_2916; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2917 = {{6'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3567 = _T_3566 + _GEN_2917; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2918 = {{7'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3568 = _T_3567 + _GEN_2918; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2919 = {{8'd0}, regs_14_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3570 = _T_3568 - _GEN_2919; // @[Conwaylife.scala 29:42]
  wire  _T_3571 = _T_3570 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3572 = _T_3570 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3573 = _T_3570 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3575 = regs_13_12 + regs_13_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2920 = {{1'd0}, regs_13_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3576 = _T_3575 + _GEN_2920; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2921 = {{2'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3577 = _T_3576 + _GEN_2921; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2922 = {{3'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3578 = _T_3577 + _GEN_2922; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2923 = {{4'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3579 = _T_3578 + _GEN_2923; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2924 = {{5'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3580 = _T_3579 + _GEN_2924; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2925 = {{6'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3581 = _T_3580 + _GEN_2925; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2926 = {{7'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3582 = _T_3581 + _GEN_2926; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2927 = {{8'd0}, regs_14_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3584 = _T_3582 - _GEN_2927; // @[Conwaylife.scala 29:42]
  wire  _T_3585 = _T_3584 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3586 = _T_3584 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3587 = _T_3584 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3589 = regs_13_13 + regs_13_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2928 = {{1'd0}, regs_13_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3590 = _T_3589 + _GEN_2928; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2929 = {{2'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3591 = _T_3590 + _GEN_2929; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2930 = {{3'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3592 = _T_3591 + _GEN_2930; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2931 = {{4'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3593 = _T_3592 + _GEN_2931; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2932 = {{5'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3594 = _T_3593 + _GEN_2932; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2933 = {{6'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3595 = _T_3594 + _GEN_2933; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2934 = {{7'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3596 = _T_3595 + _GEN_2934; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2935 = {{8'd0}, regs_14_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3598 = _T_3596 - _GEN_2935; // @[Conwaylife.scala 29:42]
  wire  _T_3599 = _T_3598 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3600 = _T_3598 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3601 = _T_3598 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3603 = regs_13_14 + regs_13_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2936 = {{1'd0}, regs_13_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3604 = _T_3603 + _GEN_2936; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2937 = {{2'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3605 = _T_3604 + _GEN_2937; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2938 = {{3'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3606 = _T_3605 + _GEN_2938; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2939 = {{4'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3607 = _T_3606 + _GEN_2939; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2940 = {{5'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3608 = _T_3607 + _GEN_2940; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2941 = {{6'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3609 = _T_3608 + _GEN_2941; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2942 = {{7'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3610 = _T_3609 + _GEN_2942; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2943 = {{8'd0}, regs_14_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3612 = _T_3610 - _GEN_2943; // @[Conwaylife.scala 29:42]
  wire  _T_3613 = _T_3612 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3614 = _T_3612 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3615 = _T_3612 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3617 = regs_14_15 + regs_14_0; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2944 = {{1'd0}, regs_14_1}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3618 = _T_3617 + _GEN_2944; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2945 = {{2'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3619 = _T_3618 + _GEN_2945; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2946 = {{3'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3620 = _T_3619 + _GEN_2946; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2947 = {{4'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3621 = _T_3620 + _GEN_2947; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2948 = {{5'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3622 = _T_3621 + _GEN_2948; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2949 = {{6'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3623 = _T_3622 + _GEN_2949; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2950 = {{7'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3624 = _T_3623 + _GEN_2950; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2951 = {{8'd0}, regs_15_0}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3626 = _T_3624 - _GEN_2951; // @[Conwaylife.scala 29:42]
  wire  _T_3627 = _T_3626 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3628 = _T_3626 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3629 = _T_3626 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3631 = regs_14_0 + regs_14_1; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2952 = {{1'd0}, regs_14_2}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3632 = _T_3631 + _GEN_2952; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2953 = {{2'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3633 = _T_3632 + _GEN_2953; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2954 = {{3'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3634 = _T_3633 + _GEN_2954; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2955 = {{4'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3635 = _T_3634 + _GEN_2955; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2956 = {{5'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3636 = _T_3635 + _GEN_2956; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2957 = {{6'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3637 = _T_3636 + _GEN_2957; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2958 = {{7'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3638 = _T_3637 + _GEN_2958; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2959 = {{8'd0}, regs_15_1}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3640 = _T_3638 - _GEN_2959; // @[Conwaylife.scala 29:42]
  wire  _T_3641 = _T_3640 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3642 = _T_3640 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3643 = _T_3640 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3645 = regs_14_1 + regs_14_2; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2960 = {{1'd0}, regs_14_3}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3646 = _T_3645 + _GEN_2960; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2961 = {{2'd0}, regs_15_1}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3647 = _T_3646 + _GEN_2961; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2962 = {{3'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3648 = _T_3647 + _GEN_2962; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2963 = {{4'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3649 = _T_3648 + _GEN_2963; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2964 = {{5'd0}, regs_0_1}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3650 = _T_3649 + _GEN_2964; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2965 = {{6'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3651 = _T_3650 + _GEN_2965; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2966 = {{7'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3652 = _T_3651 + _GEN_2966; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2967 = {{8'd0}, regs_15_2}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3654 = _T_3652 - _GEN_2967; // @[Conwaylife.scala 29:42]
  wire  _T_3655 = _T_3654 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3656 = _T_3654 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3657 = _T_3654 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3659 = regs_14_2 + regs_14_3; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2968 = {{1'd0}, regs_14_4}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3660 = _T_3659 + _GEN_2968; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2969 = {{2'd0}, regs_15_2}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3661 = _T_3660 + _GEN_2969; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2970 = {{3'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3662 = _T_3661 + _GEN_2970; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2971 = {{4'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3663 = _T_3662 + _GEN_2971; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2972 = {{5'd0}, regs_0_2}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3664 = _T_3663 + _GEN_2972; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2973 = {{6'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3665 = _T_3664 + _GEN_2973; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2974 = {{7'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3666 = _T_3665 + _GEN_2974; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2975 = {{8'd0}, regs_15_3}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3668 = _T_3666 - _GEN_2975; // @[Conwaylife.scala 29:42]
  wire  _T_3669 = _T_3668 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3670 = _T_3668 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3671 = _T_3668 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3673 = regs_14_3 + regs_14_4; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2976 = {{1'd0}, regs_14_5}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3674 = _T_3673 + _GEN_2976; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2977 = {{2'd0}, regs_15_3}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3675 = _T_3674 + _GEN_2977; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2978 = {{3'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3676 = _T_3675 + _GEN_2978; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2979 = {{4'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3677 = _T_3676 + _GEN_2979; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2980 = {{5'd0}, regs_0_3}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3678 = _T_3677 + _GEN_2980; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2981 = {{6'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3679 = _T_3678 + _GEN_2981; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2982 = {{7'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3680 = _T_3679 + _GEN_2982; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2983 = {{8'd0}, regs_15_4}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3682 = _T_3680 - _GEN_2983; // @[Conwaylife.scala 29:42]
  wire  _T_3683 = _T_3682 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3684 = _T_3682 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3685 = _T_3682 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3687 = regs_14_4 + regs_14_5; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2984 = {{1'd0}, regs_14_6}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3688 = _T_3687 + _GEN_2984; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2985 = {{2'd0}, regs_15_4}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3689 = _T_3688 + _GEN_2985; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2986 = {{3'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3690 = _T_3689 + _GEN_2986; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2987 = {{4'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3691 = _T_3690 + _GEN_2987; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2988 = {{5'd0}, regs_0_4}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3692 = _T_3691 + _GEN_2988; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2989 = {{6'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3693 = _T_3692 + _GEN_2989; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2990 = {{7'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3694 = _T_3693 + _GEN_2990; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2991 = {{8'd0}, regs_15_5}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3696 = _T_3694 - _GEN_2991; // @[Conwaylife.scala 29:42]
  wire  _T_3697 = _T_3696 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3698 = _T_3696 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3699 = _T_3696 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3701 = regs_14_5 + regs_14_6; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_2992 = {{1'd0}, regs_14_7}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3702 = _T_3701 + _GEN_2992; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_2993 = {{2'd0}, regs_15_5}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3703 = _T_3702 + _GEN_2993; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_2994 = {{3'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3704 = _T_3703 + _GEN_2994; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_2995 = {{4'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3705 = _T_3704 + _GEN_2995; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_2996 = {{5'd0}, regs_0_5}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3706 = _T_3705 + _GEN_2996; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_2997 = {{6'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3707 = _T_3706 + _GEN_2997; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_2998 = {{7'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3708 = _T_3707 + _GEN_2998; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_2999 = {{8'd0}, regs_15_6}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3710 = _T_3708 - _GEN_2999; // @[Conwaylife.scala 29:42]
  wire  _T_3711 = _T_3710 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3712 = _T_3710 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3713 = _T_3710 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3715 = regs_14_6 + regs_14_7; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3000 = {{1'd0}, regs_14_8}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3716 = _T_3715 + _GEN_3000; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3001 = {{2'd0}, regs_15_6}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3717 = _T_3716 + _GEN_3001; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3002 = {{3'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3718 = _T_3717 + _GEN_3002; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3003 = {{4'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3719 = _T_3718 + _GEN_3003; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3004 = {{5'd0}, regs_0_6}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3720 = _T_3719 + _GEN_3004; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3005 = {{6'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3721 = _T_3720 + _GEN_3005; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3006 = {{7'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3722 = _T_3721 + _GEN_3006; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3007 = {{8'd0}, regs_15_7}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3724 = _T_3722 - _GEN_3007; // @[Conwaylife.scala 29:42]
  wire  _T_3725 = _T_3724 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3726 = _T_3724 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3727 = _T_3724 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3729 = regs_14_7 + regs_14_8; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3008 = {{1'd0}, regs_14_9}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3730 = _T_3729 + _GEN_3008; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3009 = {{2'd0}, regs_15_7}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3731 = _T_3730 + _GEN_3009; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3010 = {{3'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3732 = _T_3731 + _GEN_3010; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3011 = {{4'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3733 = _T_3732 + _GEN_3011; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3012 = {{5'd0}, regs_0_7}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3734 = _T_3733 + _GEN_3012; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3013 = {{6'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3735 = _T_3734 + _GEN_3013; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3014 = {{7'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3736 = _T_3735 + _GEN_3014; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3015 = {{8'd0}, regs_15_8}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3738 = _T_3736 - _GEN_3015; // @[Conwaylife.scala 29:42]
  wire  _T_3739 = _T_3738 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3740 = _T_3738 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3741 = _T_3738 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3743 = regs_14_8 + regs_14_9; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3016 = {{1'd0}, regs_14_10}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3744 = _T_3743 + _GEN_3016; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3017 = {{2'd0}, regs_15_8}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3745 = _T_3744 + _GEN_3017; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3018 = {{3'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3746 = _T_3745 + _GEN_3018; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3019 = {{4'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3747 = _T_3746 + _GEN_3019; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3020 = {{5'd0}, regs_0_8}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3748 = _T_3747 + _GEN_3020; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3021 = {{6'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3749 = _T_3748 + _GEN_3021; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3022 = {{7'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3750 = _T_3749 + _GEN_3022; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3023 = {{8'd0}, regs_15_9}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3752 = _T_3750 - _GEN_3023; // @[Conwaylife.scala 29:42]
  wire  _T_3753 = _T_3752 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3754 = _T_3752 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3755 = _T_3752 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3757 = regs_14_9 + regs_14_10; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3024 = {{1'd0}, regs_14_11}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3758 = _T_3757 + _GEN_3024; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3025 = {{2'd0}, regs_15_9}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3759 = _T_3758 + _GEN_3025; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3026 = {{3'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3760 = _T_3759 + _GEN_3026; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3027 = {{4'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3761 = _T_3760 + _GEN_3027; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3028 = {{5'd0}, regs_0_9}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3762 = _T_3761 + _GEN_3028; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3029 = {{6'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3763 = _T_3762 + _GEN_3029; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3030 = {{7'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3764 = _T_3763 + _GEN_3030; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3031 = {{8'd0}, regs_15_10}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3766 = _T_3764 - _GEN_3031; // @[Conwaylife.scala 29:42]
  wire  _T_3767 = _T_3766 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3768 = _T_3766 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3769 = _T_3766 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3771 = regs_14_10 + regs_14_11; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3032 = {{1'd0}, regs_14_12}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3772 = _T_3771 + _GEN_3032; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3033 = {{2'd0}, regs_15_10}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3773 = _T_3772 + _GEN_3033; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3034 = {{3'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3774 = _T_3773 + _GEN_3034; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3035 = {{4'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3775 = _T_3774 + _GEN_3035; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3036 = {{5'd0}, regs_0_10}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3776 = _T_3775 + _GEN_3036; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3037 = {{6'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3777 = _T_3776 + _GEN_3037; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3038 = {{7'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3778 = _T_3777 + _GEN_3038; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3039 = {{8'd0}, regs_15_11}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3780 = _T_3778 - _GEN_3039; // @[Conwaylife.scala 29:42]
  wire  _T_3781 = _T_3780 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3782 = _T_3780 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3783 = _T_3780 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3785 = regs_14_11 + regs_14_12; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3040 = {{1'd0}, regs_14_13}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3786 = _T_3785 + _GEN_3040; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3041 = {{2'd0}, regs_15_11}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3787 = _T_3786 + _GEN_3041; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3042 = {{3'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3788 = _T_3787 + _GEN_3042; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3043 = {{4'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3789 = _T_3788 + _GEN_3043; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3044 = {{5'd0}, regs_0_11}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3790 = _T_3789 + _GEN_3044; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3045 = {{6'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3791 = _T_3790 + _GEN_3045; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3046 = {{7'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3792 = _T_3791 + _GEN_3046; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3047 = {{8'd0}, regs_15_12}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3794 = _T_3792 - _GEN_3047; // @[Conwaylife.scala 29:42]
  wire  _T_3795 = _T_3794 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3796 = _T_3794 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3797 = _T_3794 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3799 = regs_14_12 + regs_14_13; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3048 = {{1'd0}, regs_14_14}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3800 = _T_3799 + _GEN_3048; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3049 = {{2'd0}, regs_15_12}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3801 = _T_3800 + _GEN_3049; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3050 = {{3'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3802 = _T_3801 + _GEN_3050; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3051 = {{4'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3803 = _T_3802 + _GEN_3051; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3052 = {{5'd0}, regs_0_12}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3804 = _T_3803 + _GEN_3052; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3053 = {{6'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3805 = _T_3804 + _GEN_3053; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3054 = {{7'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3806 = _T_3805 + _GEN_3054; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3055 = {{8'd0}, regs_15_13}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3808 = _T_3806 - _GEN_3055; // @[Conwaylife.scala 29:42]
  wire  _T_3809 = _T_3808 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3810 = _T_3808 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3811 = _T_3808 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3813 = regs_14_13 + regs_14_14; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3056 = {{1'd0}, regs_14_15}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3814 = _T_3813 + _GEN_3056; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3057 = {{2'd0}, regs_15_13}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3815 = _T_3814 + _GEN_3057; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3058 = {{3'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3816 = _T_3815 + _GEN_3058; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3059 = {{4'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3817 = _T_3816 + _GEN_3059; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3060 = {{5'd0}, regs_0_13}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3818 = _T_3817 + _GEN_3060; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3061 = {{6'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3819 = _T_3818 + _GEN_3061; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3062 = {{7'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3820 = _T_3819 + _GEN_3062; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3063 = {{8'd0}, regs_15_14}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3822 = _T_3820 - _GEN_3063; // @[Conwaylife.scala 29:42]
  wire  _T_3823 = _T_3822 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3824 = _T_3822 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3825 = _T_3822 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [1:0] _T_3827 = regs_14_14 + regs_14_15; // @[Conwaylife.scala 29:36]
  wire [1:0] _GEN_3064 = {{1'd0}, regs_14_0}; // @[Conwaylife.scala 29:36]
  wire [2:0] _T_3828 = _T_3827 + _GEN_3064; // @[Conwaylife.scala 29:36]
  wire [2:0] _GEN_3065 = {{2'd0}, regs_15_14}; // @[Conwaylife.scala 29:36]
  wire [3:0] _T_3829 = _T_3828 + _GEN_3065; // @[Conwaylife.scala 29:36]
  wire [3:0] _GEN_3066 = {{3'd0}, regs_15_15}; // @[Conwaylife.scala 29:36]
  wire [4:0] _T_3830 = _T_3829 + _GEN_3066; // @[Conwaylife.scala 29:36]
  wire [4:0] _GEN_3067 = {{4'd0}, regs_15_0}; // @[Conwaylife.scala 29:36]
  wire [5:0] _T_3831 = _T_3830 + _GEN_3067; // @[Conwaylife.scala 29:36]
  wire [5:0] _GEN_3068 = {{5'd0}, regs_0_14}; // @[Conwaylife.scala 29:36]
  wire [6:0] _T_3832 = _T_3831 + _GEN_3068; // @[Conwaylife.scala 29:36]
  wire [6:0] _GEN_3069 = {{6'd0}, regs_0_15}; // @[Conwaylife.scala 29:36]
  wire [7:0] _T_3833 = _T_3832 + _GEN_3069; // @[Conwaylife.scala 29:36]
  wire [7:0] _GEN_3070 = {{7'd0}, regs_0_0}; // @[Conwaylife.scala 29:36]
  wire [8:0] _T_3834 = _T_3833 + _GEN_3070; // @[Conwaylife.scala 29:36]
  wire [8:0] _GEN_3071 = {{8'd0}, regs_15_15}; // @[Conwaylife.scala 29:42]
  wire [8:0] _T_3836 = _T_3834 - _GEN_3071; // @[Conwaylife.scala 29:42]
  wire  _T_3837 = _T_3836 < 9'h2; // @[Conwaylife.scala 30:16]
  wire  _T_3838 = _T_3836 == 9'h2; // @[Conwaylife.scala 32:22]
  wire  _T_3839 = _T_3836 == 9'h3; // @[Conwaylife.scala 34:22]
  wire [7:0] _T_3846 = {regs_0_7,regs_0_6,regs_0_5,regs_0_4,regs_0_3,regs_0_2,regs_0_1,regs_0_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_3854 = {regs_0_15,regs_0_14,regs_0_13,regs_0_12,regs_0_11,regs_0_10,regs_0_9,regs_0_8,_T_3846}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3861 = {regs_1_7,regs_1_6,regs_1_5,regs_1_4,regs_1_3,regs_1_2,regs_1_1,regs_1_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_3870 = {regs_1_15,regs_1_14,regs_1_13,regs_1_12,regs_1_11,regs_1_10,regs_1_9,regs_1_8,_T_3861,_T_3854}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3877 = {regs_2_7,regs_2_6,regs_2_5,regs_2_4,regs_2_3,regs_2_2,regs_2_1,regs_2_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_3885 = {regs_2_15,regs_2_14,regs_2_13,regs_2_12,regs_2_11,regs_2_10,regs_2_9,regs_2_8,_T_3877}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3892 = {regs_3_7,regs_3_6,regs_3_5,regs_3_4,regs_3_3,regs_3_2,regs_3_1,regs_3_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_3901 = {regs_3_15,regs_3_14,regs_3_13,regs_3_12,regs_3_11,regs_3_10,regs_3_9,regs_3_8,_T_3892,_T_3885}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3909 = {regs_4_7,regs_4_6,regs_4_5,regs_4_4,regs_4_3,regs_4_2,regs_4_1,regs_4_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_3917 = {regs_4_15,regs_4_14,regs_4_13,regs_4_12,regs_4_11,regs_4_10,regs_4_9,regs_4_8,_T_3909}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3924 = {regs_5_7,regs_5_6,regs_5_5,regs_5_4,regs_5_3,regs_5_2,regs_5_1,regs_5_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_3933 = {regs_5_15,regs_5_14,regs_5_13,regs_5_12,regs_5_11,regs_5_10,regs_5_9,regs_5_8,_T_3924,_T_3917}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3940 = {regs_6_7,regs_6_6,regs_6_5,regs_6_4,regs_6_3,regs_6_2,regs_6_1,regs_6_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_3948 = {regs_6_15,regs_6_14,regs_6_13,regs_6_12,regs_6_11,regs_6_10,regs_6_9,regs_6_8,_T_3940}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3955 = {regs_7_7,regs_7_6,regs_7_5,regs_7_4,regs_7_3,regs_7_2,regs_7_1,regs_7_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_3964 = {regs_7_15,regs_7_14,regs_7_13,regs_7_12,regs_7_11,regs_7_10,regs_7_9,regs_7_8,_T_3955,_T_3948}; // @[Conwaylife.scala 40:17]
  wire [127:0] _T_3966 = {_T_3964,_T_3933,_T_3901,_T_3870}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3973 = {regs_8_7,regs_8_6,regs_8_5,regs_8_4,regs_8_3,regs_8_2,regs_8_1,regs_8_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_3981 = {regs_8_15,regs_8_14,regs_8_13,regs_8_12,regs_8_11,regs_8_10,regs_8_9,regs_8_8,_T_3973}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_3988 = {regs_9_7,regs_9_6,regs_9_5,regs_9_4,regs_9_3,regs_9_2,regs_9_1,regs_9_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_3997 = {regs_9_15,regs_9_14,regs_9_13,regs_9_12,regs_9_11,regs_9_10,regs_9_9,regs_9_8,_T_3988,_T_3981}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4004 = {regs_10_7,regs_10_6,regs_10_5,regs_10_4,regs_10_3,regs_10_2,regs_10_1,regs_10_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_4012 = {regs_10_15,regs_10_14,regs_10_13,regs_10_12,regs_10_11,regs_10_10,regs_10_9,regs_10_8,_T_4004}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4019 = {regs_11_7,regs_11_6,regs_11_5,regs_11_4,regs_11_3,regs_11_2,regs_11_1,regs_11_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_4028 = {regs_11_15,regs_11_14,regs_11_13,regs_11_12,regs_11_11,regs_11_10,regs_11_9,regs_11_8,_T_4019,_T_4012}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4036 = {regs_12_7,regs_12_6,regs_12_5,regs_12_4,regs_12_3,regs_12_2,regs_12_1,regs_12_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_4044 = {regs_12_15,regs_12_14,regs_12_13,regs_12_12,regs_12_11,regs_12_10,regs_12_9,regs_12_8,_T_4036}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4051 = {regs_13_7,regs_13_6,regs_13_5,regs_13_4,regs_13_3,regs_13_2,regs_13_1,regs_13_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_4060 = {regs_13_15,regs_13_14,regs_13_13,regs_13_12,regs_13_11,regs_13_10,regs_13_9,regs_13_8,_T_4051,_T_4044}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4067 = {regs_14_7,regs_14_6,regs_14_5,regs_14_4,regs_14_3,regs_14_2,regs_14_1,regs_14_0}; // @[Conwaylife.scala 40:17]
  wire [15:0] _T_4075 = {regs_14_15,regs_14_14,regs_14_13,regs_14_12,regs_14_11,regs_14_10,regs_14_9,regs_14_8,_T_4067}; // @[Conwaylife.scala 40:17]
  wire [7:0] _T_4082 = {regs_15_7,regs_15_6,regs_15_5,regs_15_4,regs_15_3,regs_15_2,regs_15_1,regs_15_0}; // @[Conwaylife.scala 40:17]
  wire [31:0] _T_4091 = {regs_15_15,regs_15_14,regs_15_13,regs_15_12,regs_15_11,regs_15_10,regs_15_9,regs_15_8,_T_4082,_T_4075}; // @[Conwaylife.scala 40:17]
  wire [127:0] _T_4093 = {_T_4091,_T_4060,_T_4028,_T_3997}; // @[Conwaylife.scala 40:17]
  assign io_q = {_T_4093,_T_3966}; // @[Conwaylife.scala 40:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  regs_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  regs_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  regs_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  regs_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regs_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  regs_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  regs_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  regs_0_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  regs_0_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  regs_0_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  regs_0_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  regs_0_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  regs_0_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  regs_0_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  regs_0_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  regs_1_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  regs_1_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  regs_1_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  regs_1_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  regs_1_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  regs_1_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  regs_1_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  regs_1_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  regs_1_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  regs_1_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  regs_1_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  regs_1_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  regs_1_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  regs_1_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  regs_1_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  regs_1_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  regs_2_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  regs_2_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  regs_2_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  regs_2_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  regs_2_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  regs_2_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  regs_2_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  regs_2_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  regs_2_8 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  regs_2_9 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  regs_2_10 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  regs_2_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  regs_2_12 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  regs_2_13 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  regs_2_14 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  regs_2_15 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  regs_3_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  regs_3_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  regs_3_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  regs_3_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  regs_3_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  regs_3_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  regs_3_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  regs_3_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  regs_3_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  regs_3_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  regs_3_10 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  regs_3_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  regs_3_12 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  regs_3_13 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  regs_3_14 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  regs_3_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  regs_4_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  regs_4_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  regs_4_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  regs_4_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  regs_4_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  regs_4_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  regs_4_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  regs_4_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  regs_4_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  regs_4_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  regs_4_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  regs_4_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  regs_4_12 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  regs_4_13 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  regs_4_14 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  regs_4_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  regs_5_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  regs_5_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  regs_5_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  regs_5_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  regs_5_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  regs_5_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  regs_5_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  regs_5_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  regs_5_8 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  regs_5_9 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  regs_5_10 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  regs_5_11 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  regs_5_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  regs_5_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  regs_5_14 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  regs_5_15 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  regs_6_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  regs_6_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  regs_6_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  regs_6_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  regs_6_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  regs_6_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  regs_6_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  regs_6_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  regs_6_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  regs_6_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  regs_6_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  regs_6_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  regs_6_12 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  regs_6_13 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  regs_6_14 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  regs_6_15 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  regs_7_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  regs_7_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  regs_7_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  regs_7_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  regs_7_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  regs_7_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  regs_7_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  regs_7_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  regs_7_8 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  regs_7_9 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  regs_7_10 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  regs_7_11 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  regs_7_12 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  regs_7_13 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  regs_7_14 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  regs_7_15 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  regs_8_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  regs_8_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  regs_8_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  regs_8_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  regs_8_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  regs_8_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  regs_8_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  regs_8_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  regs_8_8 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  regs_8_9 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  regs_8_10 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  regs_8_11 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  regs_8_12 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  regs_8_13 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  regs_8_14 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  regs_8_15 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  regs_9_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  regs_9_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  regs_9_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  regs_9_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  regs_9_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  regs_9_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  regs_9_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  regs_9_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  regs_9_8 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  regs_9_9 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  regs_9_10 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  regs_9_11 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  regs_9_12 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  regs_9_13 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  regs_9_14 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  regs_9_15 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  regs_10_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  regs_10_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  regs_10_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  regs_10_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  regs_10_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  regs_10_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  regs_10_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  regs_10_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  regs_10_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  regs_10_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  regs_10_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  regs_10_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  regs_10_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  regs_10_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  regs_10_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  regs_10_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  regs_11_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  regs_11_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  regs_11_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  regs_11_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  regs_11_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  regs_11_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  regs_11_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  regs_11_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  regs_11_8 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  regs_11_9 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  regs_11_10 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  regs_11_11 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  regs_11_12 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  regs_11_13 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  regs_11_14 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  regs_11_15 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  regs_12_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  regs_12_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  regs_12_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  regs_12_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  regs_12_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  regs_12_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  regs_12_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  regs_12_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  regs_12_8 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  regs_12_9 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  regs_12_10 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  regs_12_11 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  regs_12_12 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  regs_12_13 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  regs_12_14 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  regs_12_15 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  regs_13_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  regs_13_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  regs_13_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  regs_13_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  regs_13_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  regs_13_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  regs_13_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  regs_13_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  regs_13_8 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  regs_13_9 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  regs_13_10 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  regs_13_11 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  regs_13_12 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  regs_13_13 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  regs_13_14 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  regs_13_15 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  regs_14_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  regs_14_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  regs_14_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  regs_14_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  regs_14_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  regs_14_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  regs_14_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  regs_14_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  regs_14_8 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  regs_14_9 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  regs_14_10 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  regs_14_11 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  regs_14_12 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  regs_14_13 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  regs_14_14 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  regs_14_15 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  regs_15_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  regs_15_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  regs_15_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  regs_15_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  regs_15_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  regs_15_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  regs_15_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  regs_15_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  regs_15_8 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  regs_15_9 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  regs_15_10 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  regs_15_11 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  regs_15_12 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  regs_15_13 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  regs_15_14 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  regs_15_15 = _RAND_255[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_load) begin
      regs_0_0 <= io_data[0];
    end else if (_T_267) begin
      regs_0_0 <= 1'h0;
    end else if (!(_T_268)) begin
      regs_0_0 <= _T_269;
    end
    if (io_load) begin
      regs_0_1 <= io_data[1];
    end else if (_T_281) begin
      regs_0_1 <= 1'h0;
    end else if (!(_T_282)) begin
      regs_0_1 <= _T_283;
    end
    if (io_load) begin
      regs_0_2 <= io_data[2];
    end else if (_T_295) begin
      regs_0_2 <= 1'h0;
    end else if (!(_T_296)) begin
      regs_0_2 <= _T_297;
    end
    if (io_load) begin
      regs_0_3 <= io_data[3];
    end else if (_T_309) begin
      regs_0_3 <= 1'h0;
    end else if (!(_T_310)) begin
      regs_0_3 <= _T_311;
    end
    if (io_load) begin
      regs_0_4 <= io_data[4];
    end else if (_T_323) begin
      regs_0_4 <= 1'h0;
    end else if (!(_T_324)) begin
      regs_0_4 <= _T_325;
    end
    if (io_load) begin
      regs_0_5 <= io_data[5];
    end else if (_T_337) begin
      regs_0_5 <= 1'h0;
    end else if (!(_T_338)) begin
      regs_0_5 <= _T_339;
    end
    if (io_load) begin
      regs_0_6 <= io_data[6];
    end else if (_T_351) begin
      regs_0_6 <= 1'h0;
    end else if (!(_T_352)) begin
      regs_0_6 <= _T_353;
    end
    if (io_load) begin
      regs_0_7 <= io_data[7];
    end else if (_T_365) begin
      regs_0_7 <= 1'h0;
    end else if (!(_T_366)) begin
      regs_0_7 <= _T_367;
    end
    if (io_load) begin
      regs_0_8 <= io_data[8];
    end else if (_T_379) begin
      regs_0_8 <= 1'h0;
    end else if (!(_T_380)) begin
      regs_0_8 <= _T_381;
    end
    if (io_load) begin
      regs_0_9 <= io_data[9];
    end else if (_T_393) begin
      regs_0_9 <= 1'h0;
    end else if (!(_T_394)) begin
      regs_0_9 <= _T_395;
    end
    if (io_load) begin
      regs_0_10 <= io_data[10];
    end else if (_T_407) begin
      regs_0_10 <= 1'h0;
    end else if (!(_T_408)) begin
      regs_0_10 <= _T_409;
    end
    if (io_load) begin
      regs_0_11 <= io_data[11];
    end else if (_T_421) begin
      regs_0_11 <= 1'h0;
    end else if (!(_T_422)) begin
      regs_0_11 <= _T_423;
    end
    if (io_load) begin
      regs_0_12 <= io_data[12];
    end else if (_T_435) begin
      regs_0_12 <= 1'h0;
    end else if (!(_T_436)) begin
      regs_0_12 <= _T_437;
    end
    if (io_load) begin
      regs_0_13 <= io_data[13];
    end else if (_T_449) begin
      regs_0_13 <= 1'h0;
    end else if (!(_T_450)) begin
      regs_0_13 <= _T_451;
    end
    if (io_load) begin
      regs_0_14 <= io_data[14];
    end else if (_T_463) begin
      regs_0_14 <= 1'h0;
    end else if (!(_T_464)) begin
      regs_0_14 <= _T_465;
    end
    if (io_load) begin
      regs_0_15 <= io_data[15];
    end else if (_T_477) begin
      regs_0_15 <= 1'h0;
    end else if (!(_T_478)) begin
      regs_0_15 <= _T_479;
    end
    if (io_load) begin
      regs_1_0 <= io_data[16];
    end else if (_T_491) begin
      regs_1_0 <= 1'h0;
    end else if (!(_T_492)) begin
      regs_1_0 <= _T_493;
    end
    if (io_load) begin
      regs_1_1 <= io_data[17];
    end else if (_T_505) begin
      regs_1_1 <= 1'h0;
    end else if (!(_T_506)) begin
      regs_1_1 <= _T_507;
    end
    if (io_load) begin
      regs_1_2 <= io_data[18];
    end else if (_T_519) begin
      regs_1_2 <= 1'h0;
    end else if (!(_T_520)) begin
      regs_1_2 <= _T_521;
    end
    if (io_load) begin
      regs_1_3 <= io_data[19];
    end else if (_T_533) begin
      regs_1_3 <= 1'h0;
    end else if (!(_T_534)) begin
      regs_1_3 <= _T_535;
    end
    if (io_load) begin
      regs_1_4 <= io_data[20];
    end else if (_T_547) begin
      regs_1_4 <= 1'h0;
    end else if (!(_T_548)) begin
      regs_1_4 <= _T_549;
    end
    if (io_load) begin
      regs_1_5 <= io_data[21];
    end else if (_T_561) begin
      regs_1_5 <= 1'h0;
    end else if (!(_T_562)) begin
      regs_1_5 <= _T_563;
    end
    if (io_load) begin
      regs_1_6 <= io_data[22];
    end else if (_T_575) begin
      regs_1_6 <= 1'h0;
    end else if (!(_T_576)) begin
      regs_1_6 <= _T_577;
    end
    if (io_load) begin
      regs_1_7 <= io_data[23];
    end else if (_T_589) begin
      regs_1_7 <= 1'h0;
    end else if (!(_T_590)) begin
      regs_1_7 <= _T_591;
    end
    if (io_load) begin
      regs_1_8 <= io_data[24];
    end else if (_T_603) begin
      regs_1_8 <= 1'h0;
    end else if (!(_T_604)) begin
      regs_1_8 <= _T_605;
    end
    if (io_load) begin
      regs_1_9 <= io_data[25];
    end else if (_T_617) begin
      regs_1_9 <= 1'h0;
    end else if (!(_T_618)) begin
      regs_1_9 <= _T_619;
    end
    if (io_load) begin
      regs_1_10 <= io_data[26];
    end else if (_T_631) begin
      regs_1_10 <= 1'h0;
    end else if (!(_T_632)) begin
      regs_1_10 <= _T_633;
    end
    if (io_load) begin
      regs_1_11 <= io_data[27];
    end else if (_T_645) begin
      regs_1_11 <= 1'h0;
    end else if (!(_T_646)) begin
      regs_1_11 <= _T_647;
    end
    if (io_load) begin
      regs_1_12 <= io_data[28];
    end else if (_T_659) begin
      regs_1_12 <= 1'h0;
    end else if (!(_T_660)) begin
      regs_1_12 <= _T_661;
    end
    if (io_load) begin
      regs_1_13 <= io_data[29];
    end else if (_T_673) begin
      regs_1_13 <= 1'h0;
    end else if (!(_T_674)) begin
      regs_1_13 <= _T_675;
    end
    if (io_load) begin
      regs_1_14 <= io_data[30];
    end else if (_T_687) begin
      regs_1_14 <= 1'h0;
    end else if (!(_T_688)) begin
      regs_1_14 <= _T_689;
    end
    if (io_load) begin
      regs_1_15 <= io_data[31];
    end else if (_T_701) begin
      regs_1_15 <= 1'h0;
    end else if (!(_T_702)) begin
      regs_1_15 <= _T_703;
    end
    if (io_load) begin
      regs_2_0 <= io_data[32];
    end else if (_T_715) begin
      regs_2_0 <= 1'h0;
    end else if (!(_T_716)) begin
      regs_2_0 <= _T_717;
    end
    if (io_load) begin
      regs_2_1 <= io_data[33];
    end else if (_T_729) begin
      regs_2_1 <= 1'h0;
    end else if (!(_T_730)) begin
      regs_2_1 <= _T_731;
    end
    if (io_load) begin
      regs_2_2 <= io_data[34];
    end else if (_T_743) begin
      regs_2_2 <= 1'h0;
    end else if (!(_T_744)) begin
      regs_2_2 <= _T_745;
    end
    if (io_load) begin
      regs_2_3 <= io_data[35];
    end else if (_T_757) begin
      regs_2_3 <= 1'h0;
    end else if (!(_T_758)) begin
      regs_2_3 <= _T_759;
    end
    if (io_load) begin
      regs_2_4 <= io_data[36];
    end else if (_T_771) begin
      regs_2_4 <= 1'h0;
    end else if (!(_T_772)) begin
      regs_2_4 <= _T_773;
    end
    if (io_load) begin
      regs_2_5 <= io_data[37];
    end else if (_T_785) begin
      regs_2_5 <= 1'h0;
    end else if (!(_T_786)) begin
      regs_2_5 <= _T_787;
    end
    if (io_load) begin
      regs_2_6 <= io_data[38];
    end else if (_T_799) begin
      regs_2_6 <= 1'h0;
    end else if (!(_T_800)) begin
      regs_2_6 <= _T_801;
    end
    if (io_load) begin
      regs_2_7 <= io_data[39];
    end else if (_T_813) begin
      regs_2_7 <= 1'h0;
    end else if (!(_T_814)) begin
      regs_2_7 <= _T_815;
    end
    if (io_load) begin
      regs_2_8 <= io_data[40];
    end else if (_T_827) begin
      regs_2_8 <= 1'h0;
    end else if (!(_T_828)) begin
      regs_2_8 <= _T_829;
    end
    if (io_load) begin
      regs_2_9 <= io_data[41];
    end else if (_T_841) begin
      regs_2_9 <= 1'h0;
    end else if (!(_T_842)) begin
      regs_2_9 <= _T_843;
    end
    if (io_load) begin
      regs_2_10 <= io_data[42];
    end else if (_T_855) begin
      regs_2_10 <= 1'h0;
    end else if (!(_T_856)) begin
      regs_2_10 <= _T_857;
    end
    if (io_load) begin
      regs_2_11 <= io_data[43];
    end else if (_T_869) begin
      regs_2_11 <= 1'h0;
    end else if (!(_T_870)) begin
      regs_2_11 <= _T_871;
    end
    if (io_load) begin
      regs_2_12 <= io_data[44];
    end else if (_T_883) begin
      regs_2_12 <= 1'h0;
    end else if (!(_T_884)) begin
      regs_2_12 <= _T_885;
    end
    if (io_load) begin
      regs_2_13 <= io_data[45];
    end else if (_T_897) begin
      regs_2_13 <= 1'h0;
    end else if (!(_T_898)) begin
      regs_2_13 <= _T_899;
    end
    if (io_load) begin
      regs_2_14 <= io_data[46];
    end else if (_T_911) begin
      regs_2_14 <= 1'h0;
    end else if (!(_T_912)) begin
      regs_2_14 <= _T_913;
    end
    if (io_load) begin
      regs_2_15 <= io_data[47];
    end else if (_T_925) begin
      regs_2_15 <= 1'h0;
    end else if (!(_T_926)) begin
      regs_2_15 <= _T_927;
    end
    if (io_load) begin
      regs_3_0 <= io_data[48];
    end else if (_T_939) begin
      regs_3_0 <= 1'h0;
    end else if (!(_T_940)) begin
      regs_3_0 <= _T_941;
    end
    if (io_load) begin
      regs_3_1 <= io_data[49];
    end else if (_T_953) begin
      regs_3_1 <= 1'h0;
    end else if (!(_T_954)) begin
      regs_3_1 <= _T_955;
    end
    if (io_load) begin
      regs_3_2 <= io_data[50];
    end else if (_T_967) begin
      regs_3_2 <= 1'h0;
    end else if (!(_T_968)) begin
      regs_3_2 <= _T_969;
    end
    if (io_load) begin
      regs_3_3 <= io_data[51];
    end else if (_T_981) begin
      regs_3_3 <= 1'h0;
    end else if (!(_T_982)) begin
      regs_3_3 <= _T_983;
    end
    if (io_load) begin
      regs_3_4 <= io_data[52];
    end else if (_T_995) begin
      regs_3_4 <= 1'h0;
    end else if (!(_T_996)) begin
      regs_3_4 <= _T_997;
    end
    if (io_load) begin
      regs_3_5 <= io_data[53];
    end else if (_T_1009) begin
      regs_3_5 <= 1'h0;
    end else if (!(_T_1010)) begin
      regs_3_5 <= _T_1011;
    end
    if (io_load) begin
      regs_3_6 <= io_data[54];
    end else if (_T_1023) begin
      regs_3_6 <= 1'h0;
    end else if (!(_T_1024)) begin
      regs_3_6 <= _T_1025;
    end
    if (io_load) begin
      regs_3_7 <= io_data[55];
    end else if (_T_1037) begin
      regs_3_7 <= 1'h0;
    end else if (!(_T_1038)) begin
      regs_3_7 <= _T_1039;
    end
    if (io_load) begin
      regs_3_8 <= io_data[56];
    end else if (_T_1051) begin
      regs_3_8 <= 1'h0;
    end else if (!(_T_1052)) begin
      regs_3_8 <= _T_1053;
    end
    if (io_load) begin
      regs_3_9 <= io_data[57];
    end else if (_T_1065) begin
      regs_3_9 <= 1'h0;
    end else if (!(_T_1066)) begin
      regs_3_9 <= _T_1067;
    end
    if (io_load) begin
      regs_3_10 <= io_data[58];
    end else if (_T_1079) begin
      regs_3_10 <= 1'h0;
    end else if (!(_T_1080)) begin
      regs_3_10 <= _T_1081;
    end
    if (io_load) begin
      regs_3_11 <= io_data[59];
    end else if (_T_1093) begin
      regs_3_11 <= 1'h0;
    end else if (!(_T_1094)) begin
      regs_3_11 <= _T_1095;
    end
    if (io_load) begin
      regs_3_12 <= io_data[60];
    end else if (_T_1107) begin
      regs_3_12 <= 1'h0;
    end else if (!(_T_1108)) begin
      regs_3_12 <= _T_1109;
    end
    if (io_load) begin
      regs_3_13 <= io_data[61];
    end else if (_T_1121) begin
      regs_3_13 <= 1'h0;
    end else if (!(_T_1122)) begin
      regs_3_13 <= _T_1123;
    end
    if (io_load) begin
      regs_3_14 <= io_data[62];
    end else if (_T_1135) begin
      regs_3_14 <= 1'h0;
    end else if (!(_T_1136)) begin
      regs_3_14 <= _T_1137;
    end
    if (io_load) begin
      regs_3_15 <= io_data[63];
    end else if (_T_1149) begin
      regs_3_15 <= 1'h0;
    end else if (!(_T_1150)) begin
      regs_3_15 <= _T_1151;
    end
    if (io_load) begin
      regs_4_0 <= io_data[64];
    end else if (_T_1163) begin
      regs_4_0 <= 1'h0;
    end else if (!(_T_1164)) begin
      regs_4_0 <= _T_1165;
    end
    if (io_load) begin
      regs_4_1 <= io_data[65];
    end else if (_T_1177) begin
      regs_4_1 <= 1'h0;
    end else if (!(_T_1178)) begin
      regs_4_1 <= _T_1179;
    end
    if (io_load) begin
      regs_4_2 <= io_data[66];
    end else if (_T_1191) begin
      regs_4_2 <= 1'h0;
    end else if (!(_T_1192)) begin
      regs_4_2 <= _T_1193;
    end
    if (io_load) begin
      regs_4_3 <= io_data[67];
    end else if (_T_1205) begin
      regs_4_3 <= 1'h0;
    end else if (!(_T_1206)) begin
      regs_4_3 <= _T_1207;
    end
    if (io_load) begin
      regs_4_4 <= io_data[68];
    end else if (_T_1219) begin
      regs_4_4 <= 1'h0;
    end else if (!(_T_1220)) begin
      regs_4_4 <= _T_1221;
    end
    if (io_load) begin
      regs_4_5 <= io_data[69];
    end else if (_T_1233) begin
      regs_4_5 <= 1'h0;
    end else if (!(_T_1234)) begin
      regs_4_5 <= _T_1235;
    end
    if (io_load) begin
      regs_4_6 <= io_data[70];
    end else if (_T_1247) begin
      regs_4_6 <= 1'h0;
    end else if (!(_T_1248)) begin
      regs_4_6 <= _T_1249;
    end
    if (io_load) begin
      regs_4_7 <= io_data[71];
    end else if (_T_1261) begin
      regs_4_7 <= 1'h0;
    end else if (!(_T_1262)) begin
      regs_4_7 <= _T_1263;
    end
    if (io_load) begin
      regs_4_8 <= io_data[72];
    end else if (_T_1275) begin
      regs_4_8 <= 1'h0;
    end else if (!(_T_1276)) begin
      regs_4_8 <= _T_1277;
    end
    if (io_load) begin
      regs_4_9 <= io_data[73];
    end else if (_T_1289) begin
      regs_4_9 <= 1'h0;
    end else if (!(_T_1290)) begin
      regs_4_9 <= _T_1291;
    end
    if (io_load) begin
      regs_4_10 <= io_data[74];
    end else if (_T_1303) begin
      regs_4_10 <= 1'h0;
    end else if (!(_T_1304)) begin
      regs_4_10 <= _T_1305;
    end
    if (io_load) begin
      regs_4_11 <= io_data[75];
    end else if (_T_1317) begin
      regs_4_11 <= 1'h0;
    end else if (!(_T_1318)) begin
      regs_4_11 <= _T_1319;
    end
    if (io_load) begin
      regs_4_12 <= io_data[76];
    end else if (_T_1331) begin
      regs_4_12 <= 1'h0;
    end else if (!(_T_1332)) begin
      regs_4_12 <= _T_1333;
    end
    if (io_load) begin
      regs_4_13 <= io_data[77];
    end else if (_T_1345) begin
      regs_4_13 <= 1'h0;
    end else if (!(_T_1346)) begin
      regs_4_13 <= _T_1347;
    end
    if (io_load) begin
      regs_4_14 <= io_data[78];
    end else if (_T_1359) begin
      regs_4_14 <= 1'h0;
    end else if (!(_T_1360)) begin
      regs_4_14 <= _T_1361;
    end
    if (io_load) begin
      regs_4_15 <= io_data[79];
    end else if (_T_1373) begin
      regs_4_15 <= 1'h0;
    end else if (!(_T_1374)) begin
      regs_4_15 <= _T_1375;
    end
    if (io_load) begin
      regs_5_0 <= io_data[80];
    end else if (_T_1387) begin
      regs_5_0 <= 1'h0;
    end else if (!(_T_1388)) begin
      regs_5_0 <= _T_1389;
    end
    if (io_load) begin
      regs_5_1 <= io_data[81];
    end else if (_T_1401) begin
      regs_5_1 <= 1'h0;
    end else if (!(_T_1402)) begin
      regs_5_1 <= _T_1403;
    end
    if (io_load) begin
      regs_5_2 <= io_data[82];
    end else if (_T_1415) begin
      regs_5_2 <= 1'h0;
    end else if (!(_T_1416)) begin
      regs_5_2 <= _T_1417;
    end
    if (io_load) begin
      regs_5_3 <= io_data[83];
    end else if (_T_1429) begin
      regs_5_3 <= 1'h0;
    end else if (!(_T_1430)) begin
      regs_5_3 <= _T_1431;
    end
    if (io_load) begin
      regs_5_4 <= io_data[84];
    end else if (_T_1443) begin
      regs_5_4 <= 1'h0;
    end else if (!(_T_1444)) begin
      regs_5_4 <= _T_1445;
    end
    if (io_load) begin
      regs_5_5 <= io_data[85];
    end else if (_T_1457) begin
      regs_5_5 <= 1'h0;
    end else if (!(_T_1458)) begin
      regs_5_5 <= _T_1459;
    end
    if (io_load) begin
      regs_5_6 <= io_data[86];
    end else if (_T_1471) begin
      regs_5_6 <= 1'h0;
    end else if (!(_T_1472)) begin
      regs_5_6 <= _T_1473;
    end
    if (io_load) begin
      regs_5_7 <= io_data[87];
    end else if (_T_1485) begin
      regs_5_7 <= 1'h0;
    end else if (!(_T_1486)) begin
      regs_5_7 <= _T_1487;
    end
    if (io_load) begin
      regs_5_8 <= io_data[88];
    end else if (_T_1499) begin
      regs_5_8 <= 1'h0;
    end else if (!(_T_1500)) begin
      regs_5_8 <= _T_1501;
    end
    if (io_load) begin
      regs_5_9 <= io_data[89];
    end else if (_T_1513) begin
      regs_5_9 <= 1'h0;
    end else if (!(_T_1514)) begin
      regs_5_9 <= _T_1515;
    end
    if (io_load) begin
      regs_5_10 <= io_data[90];
    end else if (_T_1527) begin
      regs_5_10 <= 1'h0;
    end else if (!(_T_1528)) begin
      regs_5_10 <= _T_1529;
    end
    if (io_load) begin
      regs_5_11 <= io_data[91];
    end else if (_T_1541) begin
      regs_5_11 <= 1'h0;
    end else if (!(_T_1542)) begin
      regs_5_11 <= _T_1543;
    end
    if (io_load) begin
      regs_5_12 <= io_data[92];
    end else if (_T_1555) begin
      regs_5_12 <= 1'h0;
    end else if (!(_T_1556)) begin
      regs_5_12 <= _T_1557;
    end
    if (io_load) begin
      regs_5_13 <= io_data[93];
    end else if (_T_1569) begin
      regs_5_13 <= 1'h0;
    end else if (!(_T_1570)) begin
      regs_5_13 <= _T_1571;
    end
    if (io_load) begin
      regs_5_14 <= io_data[94];
    end else if (_T_1583) begin
      regs_5_14 <= 1'h0;
    end else if (!(_T_1584)) begin
      regs_5_14 <= _T_1585;
    end
    if (io_load) begin
      regs_5_15 <= io_data[95];
    end else if (_T_1597) begin
      regs_5_15 <= 1'h0;
    end else if (!(_T_1598)) begin
      regs_5_15 <= _T_1599;
    end
    if (io_load) begin
      regs_6_0 <= io_data[96];
    end else if (_T_1611) begin
      regs_6_0 <= 1'h0;
    end else if (!(_T_1612)) begin
      regs_6_0 <= _T_1613;
    end
    if (io_load) begin
      regs_6_1 <= io_data[97];
    end else if (_T_1625) begin
      regs_6_1 <= 1'h0;
    end else if (!(_T_1626)) begin
      regs_6_1 <= _T_1627;
    end
    if (io_load) begin
      regs_6_2 <= io_data[98];
    end else if (_T_1639) begin
      regs_6_2 <= 1'h0;
    end else if (!(_T_1640)) begin
      regs_6_2 <= _T_1641;
    end
    if (io_load) begin
      regs_6_3 <= io_data[99];
    end else if (_T_1653) begin
      regs_6_3 <= 1'h0;
    end else if (!(_T_1654)) begin
      regs_6_3 <= _T_1655;
    end
    if (io_load) begin
      regs_6_4 <= io_data[100];
    end else if (_T_1667) begin
      regs_6_4 <= 1'h0;
    end else if (!(_T_1668)) begin
      regs_6_4 <= _T_1669;
    end
    if (io_load) begin
      regs_6_5 <= io_data[101];
    end else if (_T_1681) begin
      regs_6_5 <= 1'h0;
    end else if (!(_T_1682)) begin
      regs_6_5 <= _T_1683;
    end
    if (io_load) begin
      regs_6_6 <= io_data[102];
    end else if (_T_1695) begin
      regs_6_6 <= 1'h0;
    end else if (!(_T_1696)) begin
      regs_6_6 <= _T_1697;
    end
    if (io_load) begin
      regs_6_7 <= io_data[103];
    end else if (_T_1709) begin
      regs_6_7 <= 1'h0;
    end else if (!(_T_1710)) begin
      regs_6_7 <= _T_1711;
    end
    if (io_load) begin
      regs_6_8 <= io_data[104];
    end else if (_T_1723) begin
      regs_6_8 <= 1'h0;
    end else if (!(_T_1724)) begin
      regs_6_8 <= _T_1725;
    end
    if (io_load) begin
      regs_6_9 <= io_data[105];
    end else if (_T_1737) begin
      regs_6_9 <= 1'h0;
    end else if (!(_T_1738)) begin
      regs_6_9 <= _T_1739;
    end
    if (io_load) begin
      regs_6_10 <= io_data[106];
    end else if (_T_1751) begin
      regs_6_10 <= 1'h0;
    end else if (!(_T_1752)) begin
      regs_6_10 <= _T_1753;
    end
    if (io_load) begin
      regs_6_11 <= io_data[107];
    end else if (_T_1765) begin
      regs_6_11 <= 1'h0;
    end else if (!(_T_1766)) begin
      regs_6_11 <= _T_1767;
    end
    if (io_load) begin
      regs_6_12 <= io_data[108];
    end else if (_T_1779) begin
      regs_6_12 <= 1'h0;
    end else if (!(_T_1780)) begin
      regs_6_12 <= _T_1781;
    end
    if (io_load) begin
      regs_6_13 <= io_data[109];
    end else if (_T_1793) begin
      regs_6_13 <= 1'h0;
    end else if (!(_T_1794)) begin
      regs_6_13 <= _T_1795;
    end
    if (io_load) begin
      regs_6_14 <= io_data[110];
    end else if (_T_1807) begin
      regs_6_14 <= 1'h0;
    end else if (!(_T_1808)) begin
      regs_6_14 <= _T_1809;
    end
    if (io_load) begin
      regs_6_15 <= io_data[111];
    end else if (_T_1821) begin
      regs_6_15 <= 1'h0;
    end else if (!(_T_1822)) begin
      regs_6_15 <= _T_1823;
    end
    if (io_load) begin
      regs_7_0 <= io_data[112];
    end else if (_T_1835) begin
      regs_7_0 <= 1'h0;
    end else if (!(_T_1836)) begin
      regs_7_0 <= _T_1837;
    end
    if (io_load) begin
      regs_7_1 <= io_data[113];
    end else if (_T_1849) begin
      regs_7_1 <= 1'h0;
    end else if (!(_T_1850)) begin
      regs_7_1 <= _T_1851;
    end
    if (io_load) begin
      regs_7_2 <= io_data[114];
    end else if (_T_1863) begin
      regs_7_2 <= 1'h0;
    end else if (!(_T_1864)) begin
      regs_7_2 <= _T_1865;
    end
    if (io_load) begin
      regs_7_3 <= io_data[115];
    end else if (_T_1877) begin
      regs_7_3 <= 1'h0;
    end else if (!(_T_1878)) begin
      regs_7_3 <= _T_1879;
    end
    if (io_load) begin
      regs_7_4 <= io_data[116];
    end else if (_T_1891) begin
      regs_7_4 <= 1'h0;
    end else if (!(_T_1892)) begin
      regs_7_4 <= _T_1893;
    end
    if (io_load) begin
      regs_7_5 <= io_data[117];
    end else if (_T_1905) begin
      regs_7_5 <= 1'h0;
    end else if (!(_T_1906)) begin
      regs_7_5 <= _T_1907;
    end
    if (io_load) begin
      regs_7_6 <= io_data[118];
    end else if (_T_1919) begin
      regs_7_6 <= 1'h0;
    end else if (!(_T_1920)) begin
      regs_7_6 <= _T_1921;
    end
    if (io_load) begin
      regs_7_7 <= io_data[119];
    end else if (_T_1933) begin
      regs_7_7 <= 1'h0;
    end else if (!(_T_1934)) begin
      regs_7_7 <= _T_1935;
    end
    if (io_load) begin
      regs_7_8 <= io_data[120];
    end else if (_T_1947) begin
      regs_7_8 <= 1'h0;
    end else if (!(_T_1948)) begin
      regs_7_8 <= _T_1949;
    end
    if (io_load) begin
      regs_7_9 <= io_data[121];
    end else if (_T_1961) begin
      regs_7_9 <= 1'h0;
    end else if (!(_T_1962)) begin
      regs_7_9 <= _T_1963;
    end
    if (io_load) begin
      regs_7_10 <= io_data[122];
    end else if (_T_1975) begin
      regs_7_10 <= 1'h0;
    end else if (!(_T_1976)) begin
      regs_7_10 <= _T_1977;
    end
    if (io_load) begin
      regs_7_11 <= io_data[123];
    end else if (_T_1989) begin
      regs_7_11 <= 1'h0;
    end else if (!(_T_1990)) begin
      regs_7_11 <= _T_1991;
    end
    if (io_load) begin
      regs_7_12 <= io_data[124];
    end else if (_T_2003) begin
      regs_7_12 <= 1'h0;
    end else if (!(_T_2004)) begin
      regs_7_12 <= _T_2005;
    end
    if (io_load) begin
      regs_7_13 <= io_data[125];
    end else if (_T_2017) begin
      regs_7_13 <= 1'h0;
    end else if (!(_T_2018)) begin
      regs_7_13 <= _T_2019;
    end
    if (io_load) begin
      regs_7_14 <= io_data[126];
    end else if (_T_2031) begin
      regs_7_14 <= 1'h0;
    end else if (!(_T_2032)) begin
      regs_7_14 <= _T_2033;
    end
    if (io_load) begin
      regs_7_15 <= io_data[127];
    end else if (_T_2045) begin
      regs_7_15 <= 1'h0;
    end else if (!(_T_2046)) begin
      regs_7_15 <= _T_2047;
    end
    if (io_load) begin
      regs_8_0 <= io_data[128];
    end else if (_T_2059) begin
      regs_8_0 <= 1'h0;
    end else if (!(_T_2060)) begin
      regs_8_0 <= _T_2061;
    end
    if (io_load) begin
      regs_8_1 <= io_data[129];
    end else if (_T_2073) begin
      regs_8_1 <= 1'h0;
    end else if (!(_T_2074)) begin
      regs_8_1 <= _T_2075;
    end
    if (io_load) begin
      regs_8_2 <= io_data[130];
    end else if (_T_2087) begin
      regs_8_2 <= 1'h0;
    end else if (!(_T_2088)) begin
      regs_8_2 <= _T_2089;
    end
    if (io_load) begin
      regs_8_3 <= io_data[131];
    end else if (_T_2101) begin
      regs_8_3 <= 1'h0;
    end else if (!(_T_2102)) begin
      regs_8_3 <= _T_2103;
    end
    if (io_load) begin
      regs_8_4 <= io_data[132];
    end else if (_T_2115) begin
      regs_8_4 <= 1'h0;
    end else if (!(_T_2116)) begin
      regs_8_4 <= _T_2117;
    end
    if (io_load) begin
      regs_8_5 <= io_data[133];
    end else if (_T_2129) begin
      regs_8_5 <= 1'h0;
    end else if (!(_T_2130)) begin
      regs_8_5 <= _T_2131;
    end
    if (io_load) begin
      regs_8_6 <= io_data[134];
    end else if (_T_2143) begin
      regs_8_6 <= 1'h0;
    end else if (!(_T_2144)) begin
      regs_8_6 <= _T_2145;
    end
    if (io_load) begin
      regs_8_7 <= io_data[135];
    end else if (_T_2157) begin
      regs_8_7 <= 1'h0;
    end else if (!(_T_2158)) begin
      regs_8_7 <= _T_2159;
    end
    if (io_load) begin
      regs_8_8 <= io_data[136];
    end else if (_T_2171) begin
      regs_8_8 <= 1'h0;
    end else if (!(_T_2172)) begin
      regs_8_8 <= _T_2173;
    end
    if (io_load) begin
      regs_8_9 <= io_data[137];
    end else if (_T_2185) begin
      regs_8_9 <= 1'h0;
    end else if (!(_T_2186)) begin
      regs_8_9 <= _T_2187;
    end
    if (io_load) begin
      regs_8_10 <= io_data[138];
    end else if (_T_2199) begin
      regs_8_10 <= 1'h0;
    end else if (!(_T_2200)) begin
      regs_8_10 <= _T_2201;
    end
    if (io_load) begin
      regs_8_11 <= io_data[139];
    end else if (_T_2213) begin
      regs_8_11 <= 1'h0;
    end else if (!(_T_2214)) begin
      regs_8_11 <= _T_2215;
    end
    if (io_load) begin
      regs_8_12 <= io_data[140];
    end else if (_T_2227) begin
      regs_8_12 <= 1'h0;
    end else if (!(_T_2228)) begin
      regs_8_12 <= _T_2229;
    end
    if (io_load) begin
      regs_8_13 <= io_data[141];
    end else if (_T_2241) begin
      regs_8_13 <= 1'h0;
    end else if (!(_T_2242)) begin
      regs_8_13 <= _T_2243;
    end
    if (io_load) begin
      regs_8_14 <= io_data[142];
    end else if (_T_2255) begin
      regs_8_14 <= 1'h0;
    end else if (!(_T_2256)) begin
      regs_8_14 <= _T_2257;
    end
    if (io_load) begin
      regs_8_15 <= io_data[143];
    end else if (_T_2269) begin
      regs_8_15 <= 1'h0;
    end else if (!(_T_2270)) begin
      regs_8_15 <= _T_2271;
    end
    if (io_load) begin
      regs_9_0 <= io_data[144];
    end else if (_T_2283) begin
      regs_9_0 <= 1'h0;
    end else if (!(_T_2284)) begin
      regs_9_0 <= _T_2285;
    end
    if (io_load) begin
      regs_9_1 <= io_data[145];
    end else if (_T_2297) begin
      regs_9_1 <= 1'h0;
    end else if (!(_T_2298)) begin
      regs_9_1 <= _T_2299;
    end
    if (io_load) begin
      regs_9_2 <= io_data[146];
    end else if (_T_2311) begin
      regs_9_2 <= 1'h0;
    end else if (!(_T_2312)) begin
      regs_9_2 <= _T_2313;
    end
    if (io_load) begin
      regs_9_3 <= io_data[147];
    end else if (_T_2325) begin
      regs_9_3 <= 1'h0;
    end else if (!(_T_2326)) begin
      regs_9_3 <= _T_2327;
    end
    if (io_load) begin
      regs_9_4 <= io_data[148];
    end else if (_T_2339) begin
      regs_9_4 <= 1'h0;
    end else if (!(_T_2340)) begin
      regs_9_4 <= _T_2341;
    end
    if (io_load) begin
      regs_9_5 <= io_data[149];
    end else if (_T_2353) begin
      regs_9_5 <= 1'h0;
    end else if (!(_T_2354)) begin
      regs_9_5 <= _T_2355;
    end
    if (io_load) begin
      regs_9_6 <= io_data[150];
    end else if (_T_2367) begin
      regs_9_6 <= 1'h0;
    end else if (!(_T_2368)) begin
      regs_9_6 <= _T_2369;
    end
    if (io_load) begin
      regs_9_7 <= io_data[151];
    end else if (_T_2381) begin
      regs_9_7 <= 1'h0;
    end else if (!(_T_2382)) begin
      regs_9_7 <= _T_2383;
    end
    if (io_load) begin
      regs_9_8 <= io_data[152];
    end else if (_T_2395) begin
      regs_9_8 <= 1'h0;
    end else if (!(_T_2396)) begin
      regs_9_8 <= _T_2397;
    end
    if (io_load) begin
      regs_9_9 <= io_data[153];
    end else if (_T_2409) begin
      regs_9_9 <= 1'h0;
    end else if (!(_T_2410)) begin
      regs_9_9 <= _T_2411;
    end
    if (io_load) begin
      regs_9_10 <= io_data[154];
    end else if (_T_2423) begin
      regs_9_10 <= 1'h0;
    end else if (!(_T_2424)) begin
      regs_9_10 <= _T_2425;
    end
    if (io_load) begin
      regs_9_11 <= io_data[155];
    end else if (_T_2437) begin
      regs_9_11 <= 1'h0;
    end else if (!(_T_2438)) begin
      regs_9_11 <= _T_2439;
    end
    if (io_load) begin
      regs_9_12 <= io_data[156];
    end else if (_T_2451) begin
      regs_9_12 <= 1'h0;
    end else if (!(_T_2452)) begin
      regs_9_12 <= _T_2453;
    end
    if (io_load) begin
      regs_9_13 <= io_data[157];
    end else if (_T_2465) begin
      regs_9_13 <= 1'h0;
    end else if (!(_T_2466)) begin
      regs_9_13 <= _T_2467;
    end
    if (io_load) begin
      regs_9_14 <= io_data[158];
    end else if (_T_2479) begin
      regs_9_14 <= 1'h0;
    end else if (!(_T_2480)) begin
      regs_9_14 <= _T_2481;
    end
    if (io_load) begin
      regs_9_15 <= io_data[159];
    end else if (_T_2493) begin
      regs_9_15 <= 1'h0;
    end else if (!(_T_2494)) begin
      regs_9_15 <= _T_2495;
    end
    if (io_load) begin
      regs_10_0 <= io_data[160];
    end else if (_T_2507) begin
      regs_10_0 <= 1'h0;
    end else if (!(_T_2508)) begin
      regs_10_0 <= _T_2509;
    end
    if (io_load) begin
      regs_10_1 <= io_data[161];
    end else if (_T_2521) begin
      regs_10_1 <= 1'h0;
    end else if (!(_T_2522)) begin
      regs_10_1 <= _T_2523;
    end
    if (io_load) begin
      regs_10_2 <= io_data[162];
    end else if (_T_2535) begin
      regs_10_2 <= 1'h0;
    end else if (!(_T_2536)) begin
      regs_10_2 <= _T_2537;
    end
    if (io_load) begin
      regs_10_3 <= io_data[163];
    end else if (_T_2549) begin
      regs_10_3 <= 1'h0;
    end else if (!(_T_2550)) begin
      regs_10_3 <= _T_2551;
    end
    if (io_load) begin
      regs_10_4 <= io_data[164];
    end else if (_T_2563) begin
      regs_10_4 <= 1'h0;
    end else if (!(_T_2564)) begin
      regs_10_4 <= _T_2565;
    end
    if (io_load) begin
      regs_10_5 <= io_data[165];
    end else if (_T_2577) begin
      regs_10_5 <= 1'h0;
    end else if (!(_T_2578)) begin
      regs_10_5 <= _T_2579;
    end
    if (io_load) begin
      regs_10_6 <= io_data[166];
    end else if (_T_2591) begin
      regs_10_6 <= 1'h0;
    end else if (!(_T_2592)) begin
      regs_10_6 <= _T_2593;
    end
    if (io_load) begin
      regs_10_7 <= io_data[167];
    end else if (_T_2605) begin
      regs_10_7 <= 1'h0;
    end else if (!(_T_2606)) begin
      regs_10_7 <= _T_2607;
    end
    if (io_load) begin
      regs_10_8 <= io_data[168];
    end else if (_T_2619) begin
      regs_10_8 <= 1'h0;
    end else if (!(_T_2620)) begin
      regs_10_8 <= _T_2621;
    end
    if (io_load) begin
      regs_10_9 <= io_data[169];
    end else if (_T_2633) begin
      regs_10_9 <= 1'h0;
    end else if (!(_T_2634)) begin
      regs_10_9 <= _T_2635;
    end
    if (io_load) begin
      regs_10_10 <= io_data[170];
    end else if (_T_2647) begin
      regs_10_10 <= 1'h0;
    end else if (!(_T_2648)) begin
      regs_10_10 <= _T_2649;
    end
    if (io_load) begin
      regs_10_11 <= io_data[171];
    end else if (_T_2661) begin
      regs_10_11 <= 1'h0;
    end else if (!(_T_2662)) begin
      regs_10_11 <= _T_2663;
    end
    if (io_load) begin
      regs_10_12 <= io_data[172];
    end else if (_T_2675) begin
      regs_10_12 <= 1'h0;
    end else if (!(_T_2676)) begin
      regs_10_12 <= _T_2677;
    end
    if (io_load) begin
      regs_10_13 <= io_data[173];
    end else if (_T_2689) begin
      regs_10_13 <= 1'h0;
    end else if (!(_T_2690)) begin
      regs_10_13 <= _T_2691;
    end
    if (io_load) begin
      regs_10_14 <= io_data[174];
    end else if (_T_2703) begin
      regs_10_14 <= 1'h0;
    end else if (!(_T_2704)) begin
      regs_10_14 <= _T_2705;
    end
    if (io_load) begin
      regs_10_15 <= io_data[175];
    end else if (_T_2717) begin
      regs_10_15 <= 1'h0;
    end else if (!(_T_2718)) begin
      regs_10_15 <= _T_2719;
    end
    if (io_load) begin
      regs_11_0 <= io_data[176];
    end else if (_T_2731) begin
      regs_11_0 <= 1'h0;
    end else if (!(_T_2732)) begin
      regs_11_0 <= _T_2733;
    end
    if (io_load) begin
      regs_11_1 <= io_data[177];
    end else if (_T_2745) begin
      regs_11_1 <= 1'h0;
    end else if (!(_T_2746)) begin
      regs_11_1 <= _T_2747;
    end
    if (io_load) begin
      regs_11_2 <= io_data[178];
    end else if (_T_2759) begin
      regs_11_2 <= 1'h0;
    end else if (!(_T_2760)) begin
      regs_11_2 <= _T_2761;
    end
    if (io_load) begin
      regs_11_3 <= io_data[179];
    end else if (_T_2773) begin
      regs_11_3 <= 1'h0;
    end else if (!(_T_2774)) begin
      regs_11_3 <= _T_2775;
    end
    if (io_load) begin
      regs_11_4 <= io_data[180];
    end else if (_T_2787) begin
      regs_11_4 <= 1'h0;
    end else if (!(_T_2788)) begin
      regs_11_4 <= _T_2789;
    end
    if (io_load) begin
      regs_11_5 <= io_data[181];
    end else if (_T_2801) begin
      regs_11_5 <= 1'h0;
    end else if (!(_T_2802)) begin
      regs_11_5 <= _T_2803;
    end
    if (io_load) begin
      regs_11_6 <= io_data[182];
    end else if (_T_2815) begin
      regs_11_6 <= 1'h0;
    end else if (!(_T_2816)) begin
      regs_11_6 <= _T_2817;
    end
    if (io_load) begin
      regs_11_7 <= io_data[183];
    end else if (_T_2829) begin
      regs_11_7 <= 1'h0;
    end else if (!(_T_2830)) begin
      regs_11_7 <= _T_2831;
    end
    if (io_load) begin
      regs_11_8 <= io_data[184];
    end else if (_T_2843) begin
      regs_11_8 <= 1'h0;
    end else if (!(_T_2844)) begin
      regs_11_8 <= _T_2845;
    end
    if (io_load) begin
      regs_11_9 <= io_data[185];
    end else if (_T_2857) begin
      regs_11_9 <= 1'h0;
    end else if (!(_T_2858)) begin
      regs_11_9 <= _T_2859;
    end
    if (io_load) begin
      regs_11_10 <= io_data[186];
    end else if (_T_2871) begin
      regs_11_10 <= 1'h0;
    end else if (!(_T_2872)) begin
      regs_11_10 <= _T_2873;
    end
    if (io_load) begin
      regs_11_11 <= io_data[187];
    end else if (_T_2885) begin
      regs_11_11 <= 1'h0;
    end else if (!(_T_2886)) begin
      regs_11_11 <= _T_2887;
    end
    if (io_load) begin
      regs_11_12 <= io_data[188];
    end else if (_T_2899) begin
      regs_11_12 <= 1'h0;
    end else if (!(_T_2900)) begin
      regs_11_12 <= _T_2901;
    end
    if (io_load) begin
      regs_11_13 <= io_data[189];
    end else if (_T_2913) begin
      regs_11_13 <= 1'h0;
    end else if (!(_T_2914)) begin
      regs_11_13 <= _T_2915;
    end
    if (io_load) begin
      regs_11_14 <= io_data[190];
    end else if (_T_2927) begin
      regs_11_14 <= 1'h0;
    end else if (!(_T_2928)) begin
      regs_11_14 <= _T_2929;
    end
    if (io_load) begin
      regs_11_15 <= io_data[191];
    end else if (_T_2941) begin
      regs_11_15 <= 1'h0;
    end else if (!(_T_2942)) begin
      regs_11_15 <= _T_2943;
    end
    if (io_load) begin
      regs_12_0 <= io_data[192];
    end else if (_T_2955) begin
      regs_12_0 <= 1'h0;
    end else if (!(_T_2956)) begin
      regs_12_0 <= _T_2957;
    end
    if (io_load) begin
      regs_12_1 <= io_data[193];
    end else if (_T_2969) begin
      regs_12_1 <= 1'h0;
    end else if (!(_T_2970)) begin
      regs_12_1 <= _T_2971;
    end
    if (io_load) begin
      regs_12_2 <= io_data[194];
    end else if (_T_2983) begin
      regs_12_2 <= 1'h0;
    end else if (!(_T_2984)) begin
      regs_12_2 <= _T_2985;
    end
    if (io_load) begin
      regs_12_3 <= io_data[195];
    end else if (_T_2997) begin
      regs_12_3 <= 1'h0;
    end else if (!(_T_2998)) begin
      regs_12_3 <= _T_2999;
    end
    if (io_load) begin
      regs_12_4 <= io_data[196];
    end else if (_T_3011) begin
      regs_12_4 <= 1'h0;
    end else if (!(_T_3012)) begin
      regs_12_4 <= _T_3013;
    end
    if (io_load) begin
      regs_12_5 <= io_data[197];
    end else if (_T_3025) begin
      regs_12_5 <= 1'h0;
    end else if (!(_T_3026)) begin
      regs_12_5 <= _T_3027;
    end
    if (io_load) begin
      regs_12_6 <= io_data[198];
    end else if (_T_3039) begin
      regs_12_6 <= 1'h0;
    end else if (!(_T_3040)) begin
      regs_12_6 <= _T_3041;
    end
    if (io_load) begin
      regs_12_7 <= io_data[199];
    end else if (_T_3053) begin
      regs_12_7 <= 1'h0;
    end else if (!(_T_3054)) begin
      regs_12_7 <= _T_3055;
    end
    if (io_load) begin
      regs_12_8 <= io_data[200];
    end else if (_T_3067) begin
      regs_12_8 <= 1'h0;
    end else if (!(_T_3068)) begin
      regs_12_8 <= _T_3069;
    end
    if (io_load) begin
      regs_12_9 <= io_data[201];
    end else if (_T_3081) begin
      regs_12_9 <= 1'h0;
    end else if (!(_T_3082)) begin
      regs_12_9 <= _T_3083;
    end
    if (io_load) begin
      regs_12_10 <= io_data[202];
    end else if (_T_3095) begin
      regs_12_10 <= 1'h0;
    end else if (!(_T_3096)) begin
      regs_12_10 <= _T_3097;
    end
    if (io_load) begin
      regs_12_11 <= io_data[203];
    end else if (_T_3109) begin
      regs_12_11 <= 1'h0;
    end else if (!(_T_3110)) begin
      regs_12_11 <= _T_3111;
    end
    if (io_load) begin
      regs_12_12 <= io_data[204];
    end else if (_T_3123) begin
      regs_12_12 <= 1'h0;
    end else if (!(_T_3124)) begin
      regs_12_12 <= _T_3125;
    end
    if (io_load) begin
      regs_12_13 <= io_data[205];
    end else if (_T_3137) begin
      regs_12_13 <= 1'h0;
    end else if (!(_T_3138)) begin
      regs_12_13 <= _T_3139;
    end
    if (io_load) begin
      regs_12_14 <= io_data[206];
    end else if (_T_3151) begin
      regs_12_14 <= 1'h0;
    end else if (!(_T_3152)) begin
      regs_12_14 <= _T_3153;
    end
    if (io_load) begin
      regs_12_15 <= io_data[207];
    end else if (_T_3165) begin
      regs_12_15 <= 1'h0;
    end else if (!(_T_3166)) begin
      regs_12_15 <= _T_3167;
    end
    if (io_load) begin
      regs_13_0 <= io_data[208];
    end else if (_T_3179) begin
      regs_13_0 <= 1'h0;
    end else if (!(_T_3180)) begin
      regs_13_0 <= _T_3181;
    end
    if (io_load) begin
      regs_13_1 <= io_data[209];
    end else if (_T_3193) begin
      regs_13_1 <= 1'h0;
    end else if (!(_T_3194)) begin
      regs_13_1 <= _T_3195;
    end
    if (io_load) begin
      regs_13_2 <= io_data[210];
    end else if (_T_3207) begin
      regs_13_2 <= 1'h0;
    end else if (!(_T_3208)) begin
      regs_13_2 <= _T_3209;
    end
    if (io_load) begin
      regs_13_3 <= io_data[211];
    end else if (_T_3221) begin
      regs_13_3 <= 1'h0;
    end else if (!(_T_3222)) begin
      regs_13_3 <= _T_3223;
    end
    if (io_load) begin
      regs_13_4 <= io_data[212];
    end else if (_T_3235) begin
      regs_13_4 <= 1'h0;
    end else if (!(_T_3236)) begin
      regs_13_4 <= _T_3237;
    end
    if (io_load) begin
      regs_13_5 <= io_data[213];
    end else if (_T_3249) begin
      regs_13_5 <= 1'h0;
    end else if (!(_T_3250)) begin
      regs_13_5 <= _T_3251;
    end
    if (io_load) begin
      regs_13_6 <= io_data[214];
    end else if (_T_3263) begin
      regs_13_6 <= 1'h0;
    end else if (!(_T_3264)) begin
      regs_13_6 <= _T_3265;
    end
    if (io_load) begin
      regs_13_7 <= io_data[215];
    end else if (_T_3277) begin
      regs_13_7 <= 1'h0;
    end else if (!(_T_3278)) begin
      regs_13_7 <= _T_3279;
    end
    if (io_load) begin
      regs_13_8 <= io_data[216];
    end else if (_T_3291) begin
      regs_13_8 <= 1'h0;
    end else if (!(_T_3292)) begin
      regs_13_8 <= _T_3293;
    end
    if (io_load) begin
      regs_13_9 <= io_data[217];
    end else if (_T_3305) begin
      regs_13_9 <= 1'h0;
    end else if (!(_T_3306)) begin
      regs_13_9 <= _T_3307;
    end
    if (io_load) begin
      regs_13_10 <= io_data[218];
    end else if (_T_3319) begin
      regs_13_10 <= 1'h0;
    end else if (!(_T_3320)) begin
      regs_13_10 <= _T_3321;
    end
    if (io_load) begin
      regs_13_11 <= io_data[219];
    end else if (_T_3333) begin
      regs_13_11 <= 1'h0;
    end else if (!(_T_3334)) begin
      regs_13_11 <= _T_3335;
    end
    if (io_load) begin
      regs_13_12 <= io_data[220];
    end else if (_T_3347) begin
      regs_13_12 <= 1'h0;
    end else if (!(_T_3348)) begin
      regs_13_12 <= _T_3349;
    end
    if (io_load) begin
      regs_13_13 <= io_data[221];
    end else if (_T_3361) begin
      regs_13_13 <= 1'h0;
    end else if (!(_T_3362)) begin
      regs_13_13 <= _T_3363;
    end
    if (io_load) begin
      regs_13_14 <= io_data[222];
    end else if (_T_3375) begin
      regs_13_14 <= 1'h0;
    end else if (!(_T_3376)) begin
      regs_13_14 <= _T_3377;
    end
    if (io_load) begin
      regs_13_15 <= io_data[223];
    end else if (_T_3389) begin
      regs_13_15 <= 1'h0;
    end else if (!(_T_3390)) begin
      regs_13_15 <= _T_3391;
    end
    if (io_load) begin
      regs_14_0 <= io_data[224];
    end else if (_T_3403) begin
      regs_14_0 <= 1'h0;
    end else if (!(_T_3404)) begin
      regs_14_0 <= _T_3405;
    end
    if (io_load) begin
      regs_14_1 <= io_data[225];
    end else if (_T_3417) begin
      regs_14_1 <= 1'h0;
    end else if (!(_T_3418)) begin
      regs_14_1 <= _T_3419;
    end
    if (io_load) begin
      regs_14_2 <= io_data[226];
    end else if (_T_3431) begin
      regs_14_2 <= 1'h0;
    end else if (!(_T_3432)) begin
      regs_14_2 <= _T_3433;
    end
    if (io_load) begin
      regs_14_3 <= io_data[227];
    end else if (_T_3445) begin
      regs_14_3 <= 1'h0;
    end else if (!(_T_3446)) begin
      regs_14_3 <= _T_3447;
    end
    if (io_load) begin
      regs_14_4 <= io_data[228];
    end else if (_T_3459) begin
      regs_14_4 <= 1'h0;
    end else if (!(_T_3460)) begin
      regs_14_4 <= _T_3461;
    end
    if (io_load) begin
      regs_14_5 <= io_data[229];
    end else if (_T_3473) begin
      regs_14_5 <= 1'h0;
    end else if (!(_T_3474)) begin
      regs_14_5 <= _T_3475;
    end
    if (io_load) begin
      regs_14_6 <= io_data[230];
    end else if (_T_3487) begin
      regs_14_6 <= 1'h0;
    end else if (!(_T_3488)) begin
      regs_14_6 <= _T_3489;
    end
    if (io_load) begin
      regs_14_7 <= io_data[231];
    end else if (_T_3501) begin
      regs_14_7 <= 1'h0;
    end else if (!(_T_3502)) begin
      regs_14_7 <= _T_3503;
    end
    if (io_load) begin
      regs_14_8 <= io_data[232];
    end else if (_T_3515) begin
      regs_14_8 <= 1'h0;
    end else if (!(_T_3516)) begin
      regs_14_8 <= _T_3517;
    end
    if (io_load) begin
      regs_14_9 <= io_data[233];
    end else if (_T_3529) begin
      regs_14_9 <= 1'h0;
    end else if (!(_T_3530)) begin
      regs_14_9 <= _T_3531;
    end
    if (io_load) begin
      regs_14_10 <= io_data[234];
    end else if (_T_3543) begin
      regs_14_10 <= 1'h0;
    end else if (!(_T_3544)) begin
      regs_14_10 <= _T_3545;
    end
    if (io_load) begin
      regs_14_11 <= io_data[235];
    end else if (_T_3557) begin
      regs_14_11 <= 1'h0;
    end else if (!(_T_3558)) begin
      regs_14_11 <= _T_3559;
    end
    if (io_load) begin
      regs_14_12 <= io_data[236];
    end else if (_T_3571) begin
      regs_14_12 <= 1'h0;
    end else if (!(_T_3572)) begin
      regs_14_12 <= _T_3573;
    end
    if (io_load) begin
      regs_14_13 <= io_data[237];
    end else if (_T_3585) begin
      regs_14_13 <= 1'h0;
    end else if (!(_T_3586)) begin
      regs_14_13 <= _T_3587;
    end
    if (io_load) begin
      regs_14_14 <= io_data[238];
    end else if (_T_3599) begin
      regs_14_14 <= 1'h0;
    end else if (!(_T_3600)) begin
      regs_14_14 <= _T_3601;
    end
    if (io_load) begin
      regs_14_15 <= io_data[239];
    end else if (_T_3613) begin
      regs_14_15 <= 1'h0;
    end else if (!(_T_3614)) begin
      regs_14_15 <= _T_3615;
    end
    if (io_load) begin
      regs_15_0 <= io_data[240];
    end else if (_T_3627) begin
      regs_15_0 <= 1'h0;
    end else if (!(_T_3628)) begin
      regs_15_0 <= _T_3629;
    end
    if (io_load) begin
      regs_15_1 <= io_data[241];
    end else if (_T_3641) begin
      regs_15_1 <= 1'h0;
    end else if (!(_T_3642)) begin
      regs_15_1 <= _T_3643;
    end
    if (io_load) begin
      regs_15_2 <= io_data[242];
    end else if (_T_3655) begin
      regs_15_2 <= 1'h0;
    end else if (!(_T_3656)) begin
      regs_15_2 <= _T_3657;
    end
    if (io_load) begin
      regs_15_3 <= io_data[243];
    end else if (_T_3669) begin
      regs_15_3 <= 1'h0;
    end else if (!(_T_3670)) begin
      regs_15_3 <= _T_3671;
    end
    if (io_load) begin
      regs_15_4 <= io_data[244];
    end else if (_T_3683) begin
      regs_15_4 <= 1'h0;
    end else if (!(_T_3684)) begin
      regs_15_4 <= _T_3685;
    end
    if (io_load) begin
      regs_15_5 <= io_data[245];
    end else if (_T_3697) begin
      regs_15_5 <= 1'h0;
    end else if (!(_T_3698)) begin
      regs_15_5 <= _T_3699;
    end
    if (io_load) begin
      regs_15_6 <= io_data[246];
    end else if (_T_3711) begin
      regs_15_6 <= 1'h0;
    end else if (!(_T_3712)) begin
      regs_15_6 <= _T_3713;
    end
    if (io_load) begin
      regs_15_7 <= io_data[247];
    end else if (_T_3725) begin
      regs_15_7 <= 1'h0;
    end else if (!(_T_3726)) begin
      regs_15_7 <= _T_3727;
    end
    if (io_load) begin
      regs_15_8 <= io_data[248];
    end else if (_T_3739) begin
      regs_15_8 <= 1'h0;
    end else if (!(_T_3740)) begin
      regs_15_8 <= _T_3741;
    end
    if (io_load) begin
      regs_15_9 <= io_data[249];
    end else if (_T_3753) begin
      regs_15_9 <= 1'h0;
    end else if (!(_T_3754)) begin
      regs_15_9 <= _T_3755;
    end
    if (io_load) begin
      regs_15_10 <= io_data[250];
    end else if (_T_3767) begin
      regs_15_10 <= 1'h0;
    end else if (!(_T_3768)) begin
      regs_15_10 <= _T_3769;
    end
    if (io_load) begin
      regs_15_11 <= io_data[251];
    end else if (_T_3781) begin
      regs_15_11 <= 1'h0;
    end else if (!(_T_3782)) begin
      regs_15_11 <= _T_3783;
    end
    if (io_load) begin
      regs_15_12 <= io_data[252];
    end else if (_T_3795) begin
      regs_15_12 <= 1'h0;
    end else if (!(_T_3796)) begin
      regs_15_12 <= _T_3797;
    end
    if (io_load) begin
      regs_15_13 <= io_data[253];
    end else if (_T_3809) begin
      regs_15_13 <= 1'h0;
    end else if (!(_T_3810)) begin
      regs_15_13 <= _T_3811;
    end
    if (io_load) begin
      regs_15_14 <= io_data[254];
    end else if (_T_3823) begin
      regs_15_14 <= 1'h0;
    end else if (!(_T_3824)) begin
      regs_15_14 <= _T_3825;
    end
    if (io_load) begin
      regs_15_15 <= io_data[255];
    end else if (_T_3837) begin
      regs_15_15 <= 1'h0;
    end else if (!(_T_3838)) begin
      regs_15_15 <= _T_3839;
    end
  end
endmodule
